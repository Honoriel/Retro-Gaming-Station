----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 05/09/2020 09:20:59 PM
-- Design Name: 
-- Module Name: Games_Images - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use work.Defined_Values.all;


entity Games_Images is
  Port (clock, Left_button, Right_button, start_button,up_button, down_button, reset_main: in std_logic;     
        difficultyControl: in std_logic_vector(1 downto 0);  
        hSync, vSync: out std_logic;
        r, g, b: out std_logic_vector(3 downto 0));        
end Games_Images;

architecture Behavioral of Games_Images is


type success_MSG is array ( 0 to 59) of std_logic_vector( 0 to 199);
type ArrhythmiaLOGO is array (0 to 59) of std_logic_vector(0 to 299);
type ArrowGameNameMain is array (0 to 39) of std_logic_vector(0 to 159);
type Number is array (0 to 34) of std_logic_vector(0 to 89);
type Big_Number is array (0 to 79) of std_logic_vector (0 to 79);
type ArrowNotes is array (0 to 49) of std_logic_vector(0 to 49);
type ARROWMAINLOGO is array (0 to 199) of std_logic_vector(0 to 199);
type W_L_Messages is array (0 to 60) of std_logic_vector(0 to 299);
type GameStart is array (0 to 79) of std_logic_vector(0 to 399);
type InGameLogo is array (0 to 164) of std_logic_vector(0 to 199);
type PongLabel is array (0 to 63) of std_logic_vector(0 to 399);
type Main_Logos is array (0 to 299) of std_logic_vector(0 to 159);
type Selection is array (0 to 301) of std_logic_vector(0 to 161);

--Pixel Tracers
signal hPosCurrent, hPosNext: integer range 1 to H_Total;
signal vPosCurrent, vPosNext: integer range 1 to V_Total;

--RGB Signals
signal rgbCurrent, rgbNext: std_logic_vector(11 downto 0);

signal Game_Start_MessageVisible, paddleVisible,One_Three_FiveLineVisible,Two_FourLineVisible, ballVisible, paddleAIVisible,ARRHYTHMIA_GAMESTART_MESSAGEVISIBLE,ARRHYTHMIA_GAMESTART_MESSAGEVISIBLE_main, YouLoseVisible, YouWinVisible, PlayerPOINT_BITMAPVISIBLE,PlayerPOINT_BITMAP_BIGVISIBLE, AIPOINT_BITMAPVISIBLE,AIPOINT_BITMAP_BIGVISIBLE : boolean;
signal IngamelogoTopVisible,IngamelogoBottomVisible, PongNameLabelVisible, borderVisible,PongLogoVisible, ArrowLogoVisible,ArrowLogo_nameVisible, BorderLineVisible: boolean;
signal paddleCursor, paddleAICursor: integer range (H_FPorch + H_SPulse + H_BPorch + 1) to (H_Total - Width_Player):= H_FPorch + H_SPulse + H_BPorch + H_Display / 2 - (Width_Player + 1) / 2;
signal paddleLeft, paddleRight, paddleAILeft, paddleAIRight: integer range 0 to PRESCALER_PADDLE:= 0;
signal ballCursorX: integer range (H_FPorch + H_SPulse + H_BPorch + 1) to (H_Total - Ball_Size);
signal ballCursorY: integer range (V_FPorch + V_SPulse + V_BPorch + 1) to (V_Total - Ball_Size);
signal MovementCounter: integer:= 0;
signal Movement, rhythm: std_logic:= '0';
signal playingPONG, playingARROW: std_logic;
signal newGamePONG, AIWinsPONG, playerWinsPONG,AIScored, PlayerScored, newGameArrow, PlayerWonArrow, PlayerLostArrow: std_logic;
signal YouWin, YouLose: W_L_Messages;
signal GS_message: GameStart;
signal ArrowIngameLogoCircle, ArrowIngameLogoArrow : ARROWMAINLOGO;
signal UP_Arrow, Down_Arrow, Left_Arrow, Right_Arrow: ArrowNotes;
signal ArrowIngameLogoCircleVisible, ArrowIngameLogoArrowVisible, ArrowLoseVisible, ArrowWinVisible,ARRHYTHMIA_IN_GAME_Visible, UP_Coming_arrow, LEFT_Coming_arrow, RIGHT_Coming_arrow, DOWN_Coming_arrow, UP_CorrectPosition, RIGHT_CorrectPosition, LEFT_CorrectPosition, DOWN_CorrectPosition, PointVisible    : boolean :=False;
signal IngameLogoTop, IngameLogoBottom: InGameLogo;
signal PongNameLabel: PongLabel;
signal PongLogo, ArrowLogo: Main_logos;
signal AIPoint, PlayerPoint: integer range 0 to 3;
signal AIPoint_BITMAP, PlayerPoint_BITMAP: Number;
signal Borderline: Selection;
signal paddleWidth: integer:= Width_Player; 
signal WinCondition: integer range 0 to 3 ;
type screenstate is (Main,onGame1, ongame2, Game1, Game2);
signal rightbutton, leftbutton, centerbutton: integer range 0 to 35000:=0;
signal waiter: integer range 0 to 10000000:=0;
signal prev_damp: integer := 35000;
signal waitamount: integer := 10000000;
signal color_shifter: integer range 0 to 1500000:=0;
signal shifting_color: std_logic_vector := "000000000000";
signal shifting_color2: std_logic_vector := "001001001001";
signal CurrentState: screenstate := Main;
signal game_start, game_opened, Game_Opened_Arrow: std_logic:= '0';
signal UP_Current_xPOS, LEFT_Current_xPOS, RIGHT_Current_xPOS, DOWN_Current_xPOS: integer range (H_Total - H_Display + 20) to (H_Total - 30);
signal CurrentPoint: integer range 0 to 151;
signal metronome: integer range 0 to 10000000;
signal combo: std_logic := '0';
signal ArrowLogo_Name: ArrowGameNameMain;
signal ARRHYTHMIA_IN_GAME: ArrhythmiaLOGO;
signal PERFECT, GREAT, GOOD: success_MSG;
signal PerfectVisible, GreatVisible, GoodVisible: boolean := false;
signal Zero, One, Two, Three, Four, Five, Six, Seven, Eight, Nine, Ten,Eleven, Twelve, Thirteen, Fourteen, Fifteen, Sixteen, Seventeen, Eighteen, Nineteen, Twenty, Twenty_One, Twenty_Two, Twenty_Three: Number;                                       
signal Twenty_Four, Twenty_Five, Twenty_Six, Twenty_Seven, Twenty_Eight, Twenty_Nine, Thirty, Thirty_One, Thirty_Two, Thirty_Three, Thirty_Four, Thirty_Five, Thirty_Six, Thirty_Seven, Thirty_Eight, Thirty_Nine, CurrentNumber: Number;               
signal forty, forty_one, forty_two, forty_three, forty_four, forty_five, forty_six, forty_seven , forty_eight , forty_nine, fifty, fifty_one, fifty_two, fifty_three, fifty_four, fifty_five, fifty_six, fifty_seven, fifty_eight, fifty_nine: Number;                                                                                                                                                         
signal sixty, sixty_one, sixty_two, sixty_three, sixty_four, sixty_five, sixty_six, sixty_seven, sixty_eight, sixty_nine, seventy, seventy_one, seventy_two, seventy_three, seventy_four, seventy_five, seventy_six, seventy_seven, seventy_eight, seventy_nine: Number;
signal eighty, eighty_one, eighty_two, eighty_three, eighty_four, eighty_five, eighty_six, eighty_seven, eighty_eight, eighty_nine, ninety, ninety_one, ninety_two, ninety_three, ninety_four, ninety_five, ninety_six, ninety_seven, ninety_eight, ninety_nine: Number;
signal one_hundred: Number;
signal AIPoint_Bitmap_BIG, PlayerPoint_Bitmap_BIG, Zero_Big, One_big: Big_number;
signal successARROW: std_logic_vector (1 downto 0);           
signal Reaction_time, AI_Speed: integer;                                                                                                                                                                                                                                            
--Component that provides information about the balls position and game logic                                                                                                                                                                           
component PongGame is                                                                                                                                                                                                                                   
    Port (start, move, Game_on: in std_logic;                                                                                                                                                                                                           
          paddleWidth: in integer;
          WinCondition: in integer;
          AIPoint, PlayerPoint: out integer range 0 to 3;                                                                                                                                                                                                                      
          paddlePos, paddleAIPos: in integer range H_Total - H_Display + 1 to H_Total - Width_Player;                                                                                                                                                   
          xPos: out integer range H_Total - H_Display + 1 to H_Total - Ball_Size;                                                                                                                                                                       
          yPos: out integer range V_Total - V_Display + 1 to V_Total;                                                                                                                                                                                   
          newGame, play, AIWon, playerWon, AIScored, PlayerScored : out std_logic);                                                                                                                                                                                              
end component;                                                                                                                                                                                                                                          
                                                                                                                                                                                                                                                        
component ArrowGame is                                                                                                                                                                                                                                  
Port (clock, start, rhythm, Game_On, move: in std_logic;                                                                                                                                                                                                
        Up_button_Pressed, Down_button_Pressed, Left_Button_Pressed, Right_Button_Pressed: in std_logic;                                                                                                                                                
        selection_input: in std_logic_vector(1 downto 0);                                                                                                                                                                                               
        Up_xPos: out integer range (H_Total - H_Display + 20) to (H_Total - 30);                                                                                                                                                                        
        Right_xPos: out integer range (H_Total - H_Display +20) to (H_Total - 30);                                                                                                                                                                      
        Left_xPos: out integer range (H_Total - H_Display + 20) to (H_Total - 30);                                                                                                                                                                      
        Down_xPos: out integer range (H_Total - H_Display + 20) to (H_Total - 30);                                                                                                                                                                      
        newGame, play, PlayerWon, PlayerLost, on_combo: out std_logic;
        success: out std_logic_vector (1 downto 0);                                                                                                                                                                                 
        point: out integer range 0 to 151);                                                                                                                                                                                                             
end component;                                                                                                                                                                                                                                          
                                                                                                                                                                                                                                                        
                                                                                                                                                                                                                                                        
begin                                                                                                                                                                                                                                                   
    Pong: PongGame                                                                                                                                                                                                                                      
        port map (start => game_start,                                                                                                                                                                                                                  
                  move => Movement,                                                                                                                                                                                                                     
                  Game_on => Game_opened, 
                  WinCondition => WinCondition,                                                                                                                                                                                                              
                  paddleWidth => paddleWidth,                                                                                                                                                                                                           
                  paddlePos => paddleCursor,                                                                                                                                                                                                            
                  paddleAIPos => paddleAICursor,                                                                                                                                                                                                        
                  xPos => ballCursorX,                                                                                                                                                                                                                  
                  yPos => ballCursorY,                                                                                                                                                                                                                  
                  newGame => newGamePONG,                                                                                                                                                                                                               
                  play =>  playingPONG,
                  AIPoint => AIPoint,
                  PlayerPoint => PlayerPoint,                                                                                                                                                                                                                 
                  AIWon => AIWinsPONG,
                  AIScored => AIScored,
                  PlayerScored => PlayerScored,                                                                                                                                                                                                                  
                  playerWon => playerWinsPONG);                                                                                                                                                                                                         
     ArrowHero: ArrowGame                                                                                                                                                                                                                               
        port map(clock => clock,                                                                                                                                                                                                                        
                 start => game_start,                                                                                                                                                                                                                   
                 move => Movement,                                                                                                                                                                                                                      
                 rhythm => rhythm,                                                                                                                                                                                                                      
                 Game_on => Game_opened_ARROW,                                                                                                                                                                                                          
                 Up_button_Pressed => Up_button,                                                                                                                                                                                                        
                 Down_button_Pressed => Down_button,                                                                                                                                                                                                    
                 Left_Button_Pressed => Left_button,                                                                                                                                                                                                           
                 Right_Button_Pressed => Right_button,                                                                                                                                                                                                         
                 selection_input => difficultyControl,                                                                                                                                                                                                  
                 UP_xPos => UP_Current_xPOS,                                                                                                                                                                                                            
                 Right_xPos => RIGHT_Current_xPOS,                                                                                                                                                                                                      
                 Left_xPos => LEFT_Current_xPOS,                                                                                                                                                                                                        
                 Down_xPos => DOWN_Current_xPOS,                                                                                                                                                                                                        
                 point => CurrentPoint,                                                                                                                                                                                                                 
                 PlayerWon => PlayerWonArrow,                                                                                                                                                                                                           
                 PlayerLOST => PlayerLostArrow,                                                                                                                                                                                                         
                 on_combo => combo,                                                                                                                                                                                                                     
                 play => playingARROW,
                 success => successARROW,                                                                                                                                                                                                                  
                 newGame => NewGameArrow);                                                                                                                                                                                                              
                                                                                                                                                                                                                                                        
                                                                                                                                                                                                                                                        
                                                                                                                                                                                                                                                        
                                                                                                                                                                                                                                                        
                                                                                                                                                                                                                                                        
                                                                                                                                                                                                                                                        
                                                                                                                                                                                                                                                        
                                                                                                                                                                                                                                                        
process(Clock,rightbutton,leftbutton)                                                                                                                                                                                                                   
begin                                                                                                                                                                                                                                                   
if rising_edge(Clock) then                                                                                                                                                                                                                              
         if (Right_button = '1') and (Left_button= '0') then                                                                                                                                                                                                         
                            rightbutton <= rightbutton + 1;                                                                                                                                                                                             
                            leftbutton <= 0;                                                                                                                                                                                                            
                        elsif (Left_button= '1') and (Right_button = '0') then                                                                                                                                                                                       
                            leftbutton <= leftbutton + 1;                                                                                                                                                                                               
                            rightbutton <= 0;                                                                                                                                                                                                           
                        else                                                                                                                                                                                                                            
                            rightbutton <= 0;                                                                                                                                                                                                           
                            leftbutton <= 0;                                                                                                                                                                                                            
                    end if;                                                                                                                                                                                                                             
           if start_button ='1' then                                                                                                                                                                                                                    
                centerbutton <= centerbutton +1;                                                                                                                                                                                                        
           else                                                                                                                                                                                                                                         
                centerbutton <= 0;                                                                                                                                                                                                                      
           end if;                                                                                                                                                                                                                                      
          case currentstate is                                                                                                                                                                                                                          
                when Main =>                                                                                                                                                                                                                            
                    if leftbutton = prev_damp then                                                                                                                                                                                                      
                        currentstate <= onGame1;                                                                                                                                                                                                        
                    elsif rightbutton = prev_damp then                                                                                                                                                                                                  
                        currentstate <= onGame2;                                                                                                                                                                                                        
                    end if;
                when onGame1 =>
                    if centerbutton = prev_damp then
                        currentstate <= Game1;
                    elsif leftbutton = prev_damp then
                        currentstate <= onGame1;
                    elsif rightbutton = prev_damp then
                        currentstate <= onGame2;
                    end if;
                when onGame2 =>
                    if centerbutton = prev_damp then
                        currentstate <= Game2;
                    elsif leftbutton = prev_damp then
                        currentstate <= onGame1;
                    elsif rightbutton = prev_damp then
                        currentstate <= onGame2;
                    end if;
                when game1 =>
                    if game_opened ='0' then
                        waiter<= waiter + 1;
                        if waiter = waitamount then
                            game_opened<='1';
                        end if;
                    else
                        game_start <= start_button;
                    end if;
                    if reset_main ='1' then
                        currentstate <= main;
                        game_opened <='0';
                    end if;
                when game2 =>
                    if game_opened_ARROW ='0' then
                        waiter<= waiter + 1;
                        if waiter = waitamount then
                            game_opened_ARROW <='1';
                        end if;
                    else
                        game_start <= start_button;
                    end if;
                    if reset_main ='1' then
                        currentstate <= main;
                        game_opened_ARROW <='0';
                    end if;
           end case;
end if;
end process; 


    --The process involves the next state logic for the variables
    process(clock)
    begin
        if rising_edge(clock) then
            color_shifter <= color_shifter + 1;
            if color_shifter = 9999 then
                shifting_color <= std_logic_vector(unsigned(shifting_color) + 1);
                shifting_color2 <= std_logic_vector(unsigned(shifting_color2) + 1);                
            end if;
            if MovementCounter = Prescaler_Moving_Object then --Speed of the ball using a prescaler
                    Movement <= not Movement;
                    MovementCounter <= 0;
                else 
                    MovementCounter <= MovementCounter + 1;
                end if;
            if Metronome = default_rhythm then --Speed of the ball using a prescaler
                    Rhythm <= not Rhythm;
                    Metronome <= 0;
                else 
                    Metronome <= Metronome + 1;
                end if;    
                --(hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 60) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 210) and
        if currentstate = Main then
            PongLogoVisible <=(vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-150) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 150) and
                             (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + 60) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + 220) and
                                ponglogo(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-150 ))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + 60))= '0';
            ArrowLogoVisible <=(vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-150) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 150) and
                             (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 60) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 220) and
                                Arrowlogo(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-150 ))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 60))= '0';
            ArrowLogo_nameVisible <=(vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-120) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) -80) and
                                    (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 60) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 220) and
                                    ArrowLogo_Name(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-120 ))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 60))= '0';
            
            
            
            
                                                    
            hPosCurrent <= hPosNext;
            vPosCurrent <= vPosNext;
            rgbCurrent <= rgbNext;
        end if;
        if currentstate = ongame1 then
            PongLogoVisible <=(vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-150) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 150) and
                             (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + 60) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + 220) and
                                ponglogo(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-150 ))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + 60))= '0';
            ArrowLogoVisible <=(vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-150) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 150) and
                             (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 60) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 220) and
                                Arrowlogo(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-150 ))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 60))= '0';
            Borderlinevisible <= (vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-151) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 151) and
                             (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + 59) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + 221) and
                                Borderline(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-151 ))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + 59))= '0';   
             ArrowLogo_nameVisible <=(vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-120) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) -80) and
                                    (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 60) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 220) and
                                    ArrowLogo_Name(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-120 ))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 60))= '0';                              
            hPosCurrent <= hPosNext;
            vPosCurrent <= vPosNext;
            rgbCurrent <= rgbNext;
        end if;
        if currentstate = ongame2 then
            PongLogoVisible <=(vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-150) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 150) and
                             (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + 60) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + 220) and
                                ponglogo(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-150 ))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + 60))= '0';
            ArrowLogoVisible <=(vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-150) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 150) and
                             (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 60) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 220) and
                                Arrowlogo(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-150 ))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 60))= '0'; 
            Borderlinevisible <= (vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-151) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 151) and
                             (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch +(H_Display / 2)+ 59) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch+(H_Display / 2) + 221) and
                                Borderline(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-151 ))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch +(H_Display / 2)+ 59))= '0';  
             ArrowLogo_nameVisible <=(vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-120) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) -80) and
                                    (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 60) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 220) and
                                    ArrowLogo_Name(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-120 ))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 60))= '0';                                                                      
            hPosCurrent <= hPosNext;
            vPosCurrent <= vPosNext;
            rgbCurrent <= rgbNext;
        end if;
        if currentstate = game1 then
        with AIPoint select
            AIPOINT_BITMAP <= 
            Zero when 0,
            One when 1,
            two when others;
        with AIPoint select
            AIPOINT_BITMAP_BIG <= 
            Zero_BIG when 0,
            One_BIG when 1,
            ZERO_BIG when others;    
            
        
        with PlayerPoint select
            PlayerPOINT_BITMAP <= 
            Zero when 0,
            One when 1,
            two when others;
            
        with PlayerPoint select
            PlayerPOINT_BITMAP_BIG <= 
            Zero_BIG when 0,
            One_BIG when 1,
            ZERO_BIG when others;    
            
            with difficultyControl select Reaction_time <=
                        445 when "00",    
                        445 when "01",   
                        470 when "10",   
                        470 when others; 
            
            with difficultyControl select AI_SPEED <= 
                        40000 when "00",
                        40000 when "01",
                        35000 when "10",
                        35000 when others;
            with difficultyControl select WinCondition <= 
                        1 when "00",
                        2 when "01",
                        1 when "10",
                        2 when others;
            
            if playingPONG = '1' then
                if Right_button = '1' and Left_button = '0' then
                    paddleRight <= paddleRight + 1;
                    paddleLeft <= 0;
                elsif Left_button= '1' and Right_button = '0' then
                    paddleLeft <= paddleLeft + 1;
                    paddleRight <= 0;
                else 
                    paddleRight <= 0;
                    paddleLeft <= 0;
                end if;

                if paddleRight = (PRESCALER_PADDLE) and paddleCursor < H_Total - paddleWidth then
                    paddleCursor <= paddleCursor + 1;
                elsif paddleLeft = (PRESCALER_PADDLE - 5000) and paddleCursor > H_FPorch + H_SPulse + H_BPorch + 1 then
                    paddleCursor <= paddleCursor - 1;
                end if;  
                --The basic A.I algorithm with late reaction
                if (ballCursorX >= paddleAICursor) and (ballcursorY <= Reaction_Time) then --430
                    paddleAIRight <= paddleAIRight + 1;
                    paddleAILeft <= 0;
                elsif ballCursorX <= paddleAICursor and (ballcursorY <= Reaction_Time) then 
                    paddleAILeft <= paddleAILeft + 1;
                    paddleAIRight <= 0;
                else 
                    paddleAILeft <= 0;
                    paddleAIRight <= 0;
                end if;
                
                --Adjusting the position of the computer's paddle     
                if paddleAIRight = AI_SPEED and paddleAICursor < H_Total - Width_Player then
                    paddleAICursor <= paddleAICursor + 1;
                elsif paddleAILeft = AI_SPEED and paddleAICursor > H_FPorch + H_SPulse + H_BPorch + 1 then
                    paddleAICursor <= paddleAICursor - 1;
                end if;                
            else 
            
            --The initial positions of the paddles when the game stops
                paddleCursor <= H_FPorch + H_SPulse + H_BPorch + H_Display / 2 - (Width_Player + 1) / 2;
                paddleAICursor <= H_FPorch + H_SPulse + H_BPorch + H_Display / 2 - (Width_Player + 1) / 2;
            end if;
            
            hPosCurrent <= hPosNext;
            vPosCurrent <= vPosNext;
            rgbCurrent <= rgbNext;
            
   PlayerPOINT_BITMAPVISIBLE<= ( vposcurrent >=  V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 15) and ( vposcurrent <  V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 50)
                                and ( hposcurrent >= H_Total - H_display -10) and ( hposcurrent < H_Total - H_display + 80) 
                                and PlayerPoint_BITMAP(vposcurrent -( V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 15))(hposcurrent - (H_Total - H_display -10))='0' and newGamePong ='0';
   AIPOINT_BITMAPVISIBLE<= ( vposcurrent >=  V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) -50) and ( vposcurrent <  V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) -15)
                                and ( hposcurrent >= H_Total - H_display -10) and ( hposcurrent < H_Total - H_display + 80) 
                                and AIPoint_BITMAP(vposcurrent -( V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) -50))(hposcurrent - (H_Total - H_display -10))='0' and newGamePong ='0';
                                
                                
   AIPOINT_BITMAP_BIGVISIBLE<=( vposcurrent >=  V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 150) and ( vposcurrent <  V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) -70)
                              and (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 40) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 40) and
                              AIPoint_BITMAP_BIG(vposcurrent-( V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 150))(hposcurrent-( H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 40)) = '0'
                              and newGamePong ='1' and (AIscored='1' or PlayerScored ='1') and (AIWinsPong='0' and PlayerwinsPong='0');

   PlayerPOINT_BITMAP_BIGVISIBLE<=( vposcurrent >=  V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) +70) and ( vposcurrent <  V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) +150)
                              and (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 40) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 40) and
                              PlayerPoint_BITMAP_BIG(vposcurrent-( V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) +70))(hposcurrent-( H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 40)) = '0'
                              and newGamePong ='1' and (AIscored='1' or PlayerScored ='1') and (AIWinsPong='0' and PlayerwinsPong='0');
   
    YouloseVisible <= (vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 135) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 74) and
                      (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 150) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 150) and
                       YouLose(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 135))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 150)) 
                       = '0' and AIWinsPONG = '1';                  
    YouWinVisible <= (vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 135) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 74) and
                      (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 150) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 150) and
                      Youwin(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 135))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 150)) 
                      = '0' and playerWinsPONG = '1';
    Game_Start_MessageVisible <= (vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 50) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) +30) and
                      (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 200) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 200) and
                       GS_message(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 50))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 200)) 
                       = '0' and newGamePONG = '1' and ((AIWinsPONG ='0' and PlayerwinsPONG ='0' and AIScored ='0' and PlayerScored ='0')or AIwinsPONG='1' or PlayerWinsPONG ='1');
    IngamelogoTopVisible <= (vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 45) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 210) and
                   (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 100) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 100) and
                    IngamelogoTop(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 45))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 100)) 
                    = '0' and newGamePONG = '1' and ((AIWinsPONG ='0' and PlayerwinsPONG ='0' and AIScored ='0' and PlayerScored ='0')or AIwinsPONG='1' or PlayerWinsPONG ='1');
    IngamelogoBottomVisible <= (vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 45) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 210) and
                   (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 100) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 100) and
                    IngamelogoBottom(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 45))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 100)) 
                    = '0' and newGamePONG = '1' and ((AIWinsPONG ='0' and PlayerwinsPONG ='0' and AIScored ='0' and PlayerScored ='0')or AIwinsPONG='1' or PlayerWinsPONG ='1');
                                    
    PongNameLabelVisible <= (vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 150) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 86) and
                        (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 210) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 190) and
                        PongNameLabel(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 150))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 210)) 
                        = '0' and AIWinsPONG = '0' and playerWinsPONG = '0'and AIScored ='0' and PlayerScored ='0' and newGamePONG = '1';                                                                          
    paddleVisible <=    (vPosCurrent > V_Total - PADDLE_HEIGHT) and (vPosCurrent < V_Total) and (hPosCurrent >paddlecursor) and (hPosCurrent < paddlecursor + paddleWidth);
                   
    ballVisible <= ((((vPosCurrent = ballCursorY) or (vPosCurrent = ballCursorY + Ball_Size)) and (hPosCurrent > ballCursorX + 3) and (hPosCurrent <= ballCursorX + 7)) or
                   (((vPosCurrent = ballCursorY + 1) or (vPosCurrent = ballCursorY + Ball_Size - 1)) and (hPosCurrent > ballCursorX + 1) and (hPosCurrent <= ballCursorX + 9)) or
                   (((vPosCurrent = ballCursorY + 2) or (vPosCurrent = ballCursorY + Ball_Size - 2)or (vPosCurrent = ballCursorY + 3) or (vPosCurrent = ballCursorY + Ball_Size - 3)) and (hPosCurrent > ballCursorX) and (hPosCurrent <= ballCursorX + 10)) or
                   ((vPosCurrent > ballCursorY + 2) and (vPosCurrent <= ballCursorY + 7) and (hPosCurrent >= ballCursorX) and (hPosCurrent <= ballCursorX + 11))) and newGamePONG ='0' ;
    paddleAIVisible <= (vPosCurrent > V_FPorch + V_SPulse + V_BPorch  ) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch+ Paddle_HEIGHT) and (hPosCurrent >paddleAIcursor) and (hPosCurrent < paddleAIcursor + Width_Player);
                             
    borderVisible <= (vPosCurrent = V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) and newGamePONG = '0');
        end if;
        
        
        if currentstate = game2 then
     with CurrentPoint select 
     CurrentNumber <=
        Zero          when 0,
        One           when 1,
        Two           when 2,
        Three         when 3,
        Four          when 4,
        Five          when 5,
        Six           when 6,
        Seven         when 7,
        Eight         when 8,
        Nine          when 9,
        Ten           when 10,
        eleven	      when 11,
        twelve	      when 12,
        thirteen      when 13,
        fourteen      when 14,	
        fifteen	      when 15,
        sixteen	      when 16,
        seventeen     when 17,
        eighteen      when 18,	
        nineteen      when 19,	
        twenty        when 20,
        Twenty_One    when 21,
        Twenty_Two    when 22,
        Twenty_three  when 23,
        Twenty_four   when 24,
        Twenty_five   when 25,
        Twenty_six    when 26,
        Twenty_seven  when 27,
        Twenty_eight  when 28,
        Twenty_nine   when 29,
        Thirty        when 30,
        Thirty_One    when 31,
        Thirty_two    when 32,
        Thirty_three  when 33,
        Thirty_four   when 34,
        Thirty_five   when 35,
        Thirty_six    when 36,
        Thirty_seven  when 37,
        Thirty_eight  when 38,
        Thirty_nine   when 39,
        forty         when 40, 
        forty_one     when 41, 
        forty_two     when 42, 
        forty_three   when 43, 
        forty_four    when 44, 
        forty_five    when 45, 
        forty_six     when 46, 
        forty_seven   when 47, 
        forty_eight   when 48, 
        forty_nine    when 49, 
        fifty         when 50, 
        fifty_one     when 51, 
        fifty_two     when 52, 
        fifty_three   when 53, 
        fifty_four    when 54, 
        fifty_five    when 55, 
        fifty_six     when 56, 
        fifty_seven   when 57, 
        fifty_eight   when 58, 
        fifty_nine    when 59, 
        sixty         when 60, 
        sixty_one     when 61, 
        sixty_two     when 62, 
        sixty_three   when 63, 
        sixty_four    when 64, 
        sixty_five    when 65, 
        sixty_six     when 66, 
        sixty_seven   when 67, 
        sixty_eight   when 68, 
        sixty_nine    when 69, 
        seventy       when 70, 
        seventy_one   when 71, 
        seventy_two   when 72, 
        seventy_three when 73, 
        seventy_four  when 74, 
        seventy_five  when 75, 
        seventy_six   when 76, 
        seventy_seven when 77, 
        seventy_eight when 78, 
        seventy_nine  when 79, 
        eighty        when 80, 
        eighty_one    when 81, 
        eighty_two    when 82, 
        eighty_three  when 83, 
        eighty_four   when 84, 
        eighty_five   when 85, 
        eighty_six    when 86, 
        eighty_seven  when 87, 
        eighty_eight  when 88, 
        eighty_nine   when 89, 
        ninety        when 90, 
        ninety_one    when 91, 
        ninety_two    when 92, 
        ninety_three  when 93, 
        ninety_four   when 94, 
        ninety_five   when 95, 
        ninety_six    when 96, 
        ninety_seven  when 97, 
        ninety_eight  when 98, 
        ninety_nine   when 99, 
        one_hundred   when 100,
        one_hundred   when others;
        
        
     ARRHYTHMIA_GAMESTART_MESSAGEVISIBLE_Main <=(vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-100) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) -20) and
                                             (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 200) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 200) and
                                              GS_message(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 100))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 200)) 
                                              = '0' and newGameARROW = '1' and PlayerWonArrow ='0' and   PlayerLostArrow ='0';
                                              
     ARRHYTHMIA_GAMESTART_MESSAGEVISIBLE <= (vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-50) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) +30) and
                                             (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 200) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 200) and
                                              GS_message(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 50))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 200)) 
                                              = '0' and newGameARROW = '1' and (PlayerWonArrow ='1' or PlayerLostArrow ='1');   
                                                                                   
     ARRHYTHMIA_IN_GAME_Visible <= (vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) -200) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-140) and 
                                     (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 150) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 150) and
                                     ARRHYTHMIA_IN_GAME(vPosCurrent -( V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 200))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 150))='0' 
                                     and newGameArrow ='1' and PlayerWonArrow ='0' and   PlayerLostArrow ='0';
     
     
     ArrowIngameLogoCircleVisible <= (vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) ) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 200) and 
                                     (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 100) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 100) and
                                     ArrowIngameLogoCircle(vPosCurrent -( V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 100))='0' 
                                     and newGameArrow ='1' and PlayerWonArrow ='0' and   PlayerLostArrow ='0';
                                                                
     
     ArrowIngameLogoArrowVisible <=  (vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) ) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 200) and 
                                     (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 100) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 100) and
                                     ArrowIngameLogoArrow(vPosCurrent -( V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 100))='0' 
                                     and newGameArrow ='1' and PlayerWonArrow ='0' and   PlayerLostArrow ='0';
                                     
     One_Three_FiveLineVisible <=  (hposcurrent > H_Total - H_Display + 60) and (hposcurrent < H_Total -25) and ((Vposcurrent = V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 210) or (Vposcurrent = V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 50)
                                     or (Vposcurrent = V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 110))and newGameArrow ='0' ;
     Two_FourLineVisible <= (hposcurrent >H_Total - H_Display + 60) and (hposcurrent < H_Total -25) and ((Vposcurrent = V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 126)or (Vposcurrent = V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 26))and newGameArrow ='0' ;
                                                                
     ArrowWinVisible <=(vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 135) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 74) and
                      (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 150) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 150) and
                       YouWin(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 135))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 150)) 
                       = '0' and PlayerWonArrow = '1';
    
                                  
     ArrowLoseVisible <=(vPosCurrent >= V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 135) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 74) and
                      (hPosCurrent >= H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 150) and (hPosCurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) + 150) and
                       YouLose(vPosCurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 135))(hPosCurrent - (H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) - 150)) 
                       = '0' and PlayerLostArrow = '1';
     
     UP_Coming_arrow <= (Hposcurrent > UP_Current_xPOS )and (Hposcurrent < UP_Current_xPOS +50) and (vPosCurrent > V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 195) and(vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 145) and
                        UP_Arrow(vposcurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 195))(Hposcurrent - up_Current_xPos) ='0'  and newGameArrow ='0' ;
                        
     LEFT_Coming_arrow <= (Hposcurrent > LEFT_Current_xPOS )and (Hposcurrent < LEFT_Current_xPOS +50) and (vPosCurrent > V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 115) and(vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) -65) and 
                           LEFT_Arrow(vposcurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 115))(Hposcurrent - left_Current_xPos) ='0'  and newGameArrow ='0' ;
          
     RIGHT_Coming_arrow <= (Hposcurrent > RIGHT_Current_xPOS )and (Hposcurrent < RIGHT_Current_xPOS +50)and (vPosCurrent > V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 35) and(vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 15) and
                            RIGHT_Arrow(vposcurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-35))(Hposcurrent - right_Current_xPos) ='0'  and newGameArrow ='0' ;

     DOWN_Coming_arrow <= (Hposcurrent > DOWN_Current_xPOS )and (Hposcurrent < DOWN_Current_xPOS +50)and (vPosCurrent > V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 45) and(vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 95) and 
                            DOWN_Arrow(vposcurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 45))(Hposcurrent - down_Current_xPos) ='0'  and newGameArrow ='0' ;

     
     Up_CorrectPosition <= (hposcurrent < H_Total - H_Display + 83) and (hposcurrent > H_Total - H_Display + 33)and (vPosCurrent > V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 195) and(vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 145) and
                            UP_Arrow(vposcurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 195))(Hposcurrent - (H_Total - H_Display + 33)) ='0'  and newGameArrow ='0' ; 
     
     
     LEFT_CorrectPosition <=  (hposcurrent < H_Total - H_Display + 83) and (hposcurrent > H_Total - H_Display + 33)and (vPosCurrent > V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 115) and(vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 65) and                                    
                               LEFT_Arrow(vposcurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) - 115))(Hposcurrent - (H_Total - H_Display + 33)) ='0'  and newGameArrow ='0' ;                                                                                                    
     
     RIGHT_CorrectPosition <= (hposcurrent < H_Total - H_Display + 83) and (hposcurrent > H_Total - H_Display + 33)and (vPosCurrent > V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-35 ) and(vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 15) and                
                                 RIGHT_Arrow(vposcurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)-35))(Hposcurrent - (H_Total - H_Display + 33)) ='0'  and newGameArrow ='0' ; 
                                 
     DOWN_CorrectPosition <= (hposcurrent < H_Total - H_Display + 83) and (hposcurrent > H_Total - H_Display + 33)and (vPosCurrent > V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 45) and(vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 95) and                
                                DOWN_Arrow(vposcurrent - (V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) +45))(Hposcurrent - (H_Total - H_Display + 33)) ='0'  and newGameArrow ='0' ;                                                                                                                                
                                                                                                                                    
     PointVisible <= (hposcurrent < H_Total - H_Display + 120) and (hposcurrent > H_Total - H_Display + 30)and (vPosCurrent > V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 160) and (vPosCurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 195) 
                    and CurrentNumber(vposcurrent -(V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 160))(hposcurrent-(H_Total - H_Display + 30))='0' and (newGameArrow ='0' or PlayerWonArrow = '1' or PlayerLostArrow = '1');
     
     PerfectVisible<= (vposcurrent >  V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 60) and (vposcurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)+120)
                      and (hposcurrent > H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) -100) and ( hposcurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2)+100)
                      and PERFECT(vposcurrent -(V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 60))(hposcurrent-(H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) -100))='0' and successARROW ="11"  and PlayerWonArrow = '1';
     
     
     GreatVisible  <=(vposcurrent >  V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 60) and (vposcurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)+120)
                      and (hposcurrent > H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) -100) and ( hposcurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2)+100)
                      and Great(vposcurrent -(V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 60))(hposcurrent-(H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) -100))='0' and successARROW ="10"  and PlayerWonArrow = '1';
     
     
     GoodVisible   <=(vposcurrent >  V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 60) and (vposcurrent < V_FPorch + V_SPulse + V_BPorch + (V_Display / 2)+120)
                      and (hposcurrent > H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) -100) and ( hposcurrent < H_FPorch + H_SPulse + H_BPorch + (H_Display / 2)+100)
                      and GOOD(vposcurrent -(V_FPorch + V_SPulse + V_BPorch + (V_Display / 2) + 60))(hposcurrent-(H_FPorch + H_SPulse + H_BPorch + (H_Display / 2) -100))='0' and successARROW ="01"  and PlayerWonArrow = '1';
     
     
            hPosCurrent <= hPosNext;
            vPosCurrent <= vPosNext;
            rgbCurrent <= rgbNext;
        
        end if;
        end if;
    end process;

    --Scanning the Pixels with predefined values:
    hPosNext <= hPosCurrent + 1 when hPosCurrent < H_Total else 1;
    vPosNext <= vPosCurrent + 1 when hPosCurrent = H_Total and vPosCurrent < V_Total else
                1 when hPosCurrent = H_Total and vPosCurrent = V_Total else vPosCurrent;
        
        
        
        -- color assignments to display images
        rgbNext <= "111111111111"  when PonglogoVisible or PLayerPoint_bitmapvisible or AIPoint_bitmapvisible  or ARRHYTHMIA_GAMESTART_MESSAGEVISIBLE or ARRHYTHMIA_GAMESTART_MESSAGEVISIBLE_main  or PlayerPOINT_BITMAP_BIGVISIBLE or AIPOINT_BITMAP_BIGVISIBLE or ArrowLogo_nameVisible or ARRHYTHMIA_IN_GAME_Visible else
                   "001001110111"  when BorderlineVisible else 
                   shifting_color  when Arrowlogovisible or One_Three_FiveLineVisible  else --"111100001111"
                   shifting_color2 when Two_FourLineVisible or PerfectVisible else
                   "111111111111"  when paddleVisible else
                   "111111111111"  when Game_Start_MessageVisible else
                   "111011101110"  when ballVisible else                     
                   "111111111111"  when borderVisible else
                   "111100000000"  when paddleAIVisible else 
                   "000011111111"  when YouWinVisible else
                   "111100000000"  when YouLoseVisible else
                   "111100000000"  when ArrowLoseVisible else
                   "000011111111"  when ArrowWinVisible or GreatVisible else
                   "111111111111"  when PongNameLabelVisible or GoodVisible else
                   "111111111111"  when IngamelogoTopVisible else
                   "111111110111"  when IngamelogoBottomVisible else
                   "010100000110"  when ArrowIngameLogoCircleVisible else
                   shifting_color  when ArrowIngameLogoArrowVisible else
                   "111111111111"  when UP_Coming_arrow or LEFT_Coming_arrow or RIGHT_Coming_arrow or DOWN_Coming_arrow or Pointvisible else
                   "101010101010"  when Up_CorrectPosition or RIght_CorrectPosition or LEFT_CorrectPosition or DOWN_CorrectPosition  else
                   "000000000000";    
                   
    --Updating rgb and hsync, vsync 
    hSync <= '0' when (hPosCurrent > H_FPorch) and (hPosCurrent < H_FPorch + H_SPulse + 1) else '1';
    vSync <= '0' when (vPosCurrent > V_FPorch) and (vPosCurrent < V_FPorch + V_SPulse + 1) else '1';
    r <= rgbCurrent(11 downto 8);
    g <= rgbCurrent(7 downto 4);
    b <= rgbCurrent(3 downto 0);    

   YouWin<=("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
            "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
            "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
            "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111",
            "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111",
            "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111",
            "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000111111",
            "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000011",
            "111111111111111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000011",
            "110000000000000000000000000000001111111111110000000000000000000000000011111111110000000000000001111000000000000000111111111111111111111111111111111000000000000000111000000000000000111111111111000000000000000000000000001111111111000000000000000111000000000000000111111111111110000011111111000000000011",
            "110000000000000000000000000000001111111111110000000000000000000000000011111111110000000000000001111000000000000000111111111111111111111111111111111000000000000000111000000000000000111111111111000000000000000000000000001111111111000000000000000111000000000000000111111111111110000011111111000000000011",
            "110000000000000000000000000000001111111111110000000000000000000000000011111111110000000000000001111000000000000000111111111111111111111111111111111000000000000000111000000000000000111111111111000000000000000000000000001111111111000000000000000111000000000000000111111111111110000011111111000000000011",
            "110000000000000000000000000000001111111111110000000000000000000000000011111111110000000000000001111000000000000000111111111111111111111111111111111000000000000000111000000000000000111111111111000000000000000000000000001111111111000000000000000111000000000000000111111111111110000011111111000000000011",
            "110000000000000000000000000000001111111100000001111111111111111111000000011111110000000000000000111000000000000000111111111111111111111111111111111000000000000000111000000000000000111111111111000000000000000000000000001111111111000000000000000111000000000000000111111111111110000011111111000000000011",
            "110000111111100000001111111100000000111100000001111111111111111111000000011111110000111111110000000000011111110000000111111111111111111111111111111000011111110000000000001111111000000011110000000011111111111111111100000001111111000011111110000000000001111110000000011111111110000011111111000000000011",
            "110000111111100000001111111100000001111100000001111111111111111111000000011111110000111111110000000000011111110000000111111111111111111111111111111000011111110000000000011111111000000011110000000111111111111111111100000001111111000011111110000000000011111111000000011111111110000011111111000000000011",
            "110000111111100000001111111100000001111100000001111111111111111111000000011111110000111111110000000000011111110000000111111111111111111111111111111000011111110000000000011111111000000011110000000111111111111111111100000001111111000011111110000000000011111111000000011111111110000011111111000000000011",
            "110000111111100000001111111100000001111100000001111111111111111111000000001111110000111111110000000000011111110000000111111111111111111111111111111000011111110000000000011111111000000011110000000111111111111111111100000001111111000011111110000000000011111111000000011111111110000011111111000000000011",
            "110000111111100000001111111100000001111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111110000000000011111111000000011110000000111111111111111111100000001111111000011111110000000000011111111000000011111111110000011111111000000000011",
            "110000111111100000001111111100000001111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111110000000000011111111000000011110000111111100000000000111111110000000111000011111111111000000011111111000000011111111110000011111111000000000011",
            "110000111111100000001111111100000001111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111110000000000011111111000000011110000111111100000000000111111110000000111000011111111111000000011111111000000011111111110000011111111000000000011",
            "110000111111100000001111111100000001111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111110000000000011111111000000011110000111111100000000000111111110000000111000011111111111000000011111111000000011111111110000011111111000000000011",
            "110000111111100000001111111100000001111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111110000000000011111111000000011110000111111100000000000111111110000000111000011111111111000000011111111000000011111111110000011111111000000000011",
            "110000111111100000001111111100000001111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111110000000000011111111000000011110000111111100000000000111111110000000111000011111111111111000011111111000000011111111110000011111111000000000011",
            "110000111111100000001111111100000001111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111110000000000011111111000000011110000111111100000000000111111110000000111000011111111111111000011111111000000011111111110000011111111000000000011",
            "110000111111100000001111111100000001111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111110000000000011111111000000011110000111111100000000000111111110000000111000011111111111111000011111111000000011111111110000011111000000000000011",
            "110000111111100000001111111100000001111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111110000000000011111111000000011110000111111100000000000111111110000000111000011111111111111000011111111000000011111111110000011111000000000000011",
            "110000000111111111111111000000000001111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111110000000000011111111000000011110000111111100000000000111111110000000111000011111111111111000011111111000000011111111110000011111000000000000011",
            "110000000111111111111111000000000001111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111110000111000011111111000000011110000111111100000000000111111110000000111000011111110000111111111111111000000011111111110000011111000000000000011",
            "110000000111111111111111000000000001111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111110000111000011111111000000011110000111111100000000000111111110000000111000011111110000111111111111111000000011111111110000011111000000000000011",
            "110000000111111111111111000000000001111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111110000111000011111111000000011110000111111100000000000111111110000000111000011111110000111111111111111000000011111111110000011111000000000000011",
            "110000000111111111111111000000000001111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111110000111000011111111000000011110000111111100000000000111111110000000111000011111110000111111111111111000000011111111110000011111000000000000011",
            "111111000000011111110000000000000001111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111111111111111111111111000000011110000111111100000000000111111110000000111000011111110000111111111111111000000011111111110000011111000000000000011",
            "111111000000011111110000000000000001111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111111111111111111111111000000011110000111111100000000000111111110000000111000011111110000000111111111111000000011111111110000011110000000000000011",
            "111111000000011111110000000000000001111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111111111111111111111111000000011110000111111100000000000111111110000000111000011111110000000111111111111000000011111111110000011110000000000000011",
            "111111000000011111110000000000000000111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111111111111111111111111000000011110000111111100000000000111111110000000111000011111110000000111111111111000000011111111110000011110000000000111111",
            "111111000000011111110000000000000001111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111111111111111111111111000000011110000111111100000000000111111110000000111000011111110000000111111111111000000011111111110000011110000000000111111",
            "111111111000011111110000000000001111111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111111111000111111111111000000011110000111111100000000000111111110000000111000011111110000000111111111111000000011111111110000000000000000000111111",
            "111111111000011111110000000000001111111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111111111000111111111111000000011110000111111100000000000111111110000000111000011111110000000000011111111000000011111111110000000000000000000111111",
            "111111111000011111110000000000001111111100001111111000000000001111111100000001110000111111110000000000011111110000000111111111111111111111111111111000011111111111000111111111111000000011110000111111100000000000111111110000000111000011111110000000000011111111000000011111111110000000000000000000111111",
            "111111111000011111110000000000001111111100000001111111111111111111000000000001110000111111110000000000011111110000000111111111111111111111111111111000011111111111000111111111111000000011110000111111100000000000111111110000000111000011111110000000000011111111000000011111111110000000000000000000111111",
            "111111111000011111110000000011111111111100000001111111111111111111000000000001110000000011111111111111111100000000000111111111111111111111111111111000011111111111000111111111111000000011110000111111110000000000111111110000000111000011111110000000000011111111000000011111111110000011110000000000111111",
            "111111111000011111110000000011111111111100000001111111111111111111000000000001110000000011111111111111111100000000000111111111111111111111111111111000011111110000000000011111111000000011110000000111111111111111111100000000000111000011111110000000000011111111000000011111111110000011110000000000111111",
            "111111111000011111110000000011111111111100000001111111111111111111000000000001110000000011111111111111111100000000000111111111111111111111111111111000011111110000000000011111111000000011110000000111111111111111111100000000000111000011111110000000000011111111000000011111111110000011110000000000111111",
            "111111111000011111110000000011111111111100000001111111111111111111000000000001110000000011111111111111111100000000000111111111111111111111111111111000011111110000000000011111111000000011110000000111111111111111111100000000000111000011111110000000000011111111000000011111111110000011110000000000111111",
            "111111111000011111110000000011111111111100000000111111111111111111000000000001110000000011111111111111111100000000000111111111111111111111111111111000011111110000000000011111111000000011110000000111111111111111111100000000000111000011111110000000000011111111000000011111111110000011110000000000111111",
            "111111111000000000000000000011111111111111110000000000000000000000000000000001111111000000000000000000000000000000000111111111111111111111111111111000011111110000000000011111111000000011110000000111111111111111111100000000000111000011111110000000000001111110000000011111111110000011110000000000111111",
            "111111111000000000000000000011111111111111110000000000000000000000000000000001111111000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000011111111000000000000000000000000000000000111000000000000000000000000000000000000011111111110000011110000000000111111",
            "111111111000000000000000000011111111111111110000000000000000000000000000000001111111000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000011111111000000000000000000000000000000000111000000000000000000000000000000000000011111111110000000000000000000111111",
            "111111111000000000000000000011111111111111110000000000000000000000000000000001111111000000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000011111111000000000000000000000000000000000111000000000000000000000000000000000000011111111110000000000000000000111111",
            "111111111100000000000000000011111111111111111110000000000000000000000000011111111111100000000000000000000000000000000111111111111111111111111111111000000000000000000000000000000000000011111111000000000000000000000000000000000111000000000000000000000000000000000000011111111110000000000000000000111111",
            "111111111111100000000000000011111111111111111110000000000000000000000000011111111111111100000000000000000000000000111111111111111111111111111111111111100000000000000011100000000000000011111111111000000000000000000000000000111111111100000000000000111100000000000000011111111110000000000000000000111111",
            "111111111111100000000000000011111111111111111110000000000000000000000000011111111111111100000000000000000000000000111111111111111111111111111111111111100000000000000111100000000000000011111111111000000000000000000000000001111111111100000000000000111100000000000000011111111110000000000000000000111111",
            "111111111111100000000000000011111111111111111110000000000000000000000000011111111111111100000000000000000000000000111111111111111111111111111111111111100000000000000111100000000000000011111111111000000000000000000000000001111111111100000000000000111100000000000000011111111111111100000000000000111111",
            "111111111111100000000000000011111111111111111111000000000000000000000000011111111111111100000000000000000000000000111111111111111111111111111111111111100000000000000111100000000000000011111111111000000000000000000000000001111111111100000000000000111100000000000000011111111111111100000000000000111111",
            "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111100000000000000011111111111000000000000000000000000001111111111100000000000000111100000000000000011111111111111100000000000000111111",
            "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111",
            "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111",
            "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111",
            "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
            "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");
            
    YouLose <=("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
               "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
               "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111", 
               "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111", 
               "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111", 
               "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111", 
               "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000011111", 
               "110000000000000000000000000000111111111110000000000000000000000000111111111000000000000001110000000000000011111111111111111111111000000000000001111111111111111111111110000000000000000000000000111111111111100000000000000000000000011111111110000000000000000000000000000111111111100000000000000000000011", 
               "110000000000000000000000000000111111111110000000000000000000000001111111111000000000000001110000000000000011111111111111111111111000000000000001111111111111111111111110000000000000000000000000111111111111100000000000000000000000011111111110000000000000000000000000000111111111100000000000000000000011", 
               "110000000000000000000000000000111111111110000000000000000000000001111111111000000000000001110000000000000011111111111111111111111000000000000001111111111111111111111110000000000000000000000000111111111111100000000000000000000000011111111110000000000000000000000000000111111111100001111111100000000011", 
               "110000000000000000000000000000111111111110000000000000000000000001111111111000000000000001110000000000000011111111111111111111111000000000000001111111111111111111111110000000000000000000000000111111111111100000000000000000000000011111111110000000000000000000000000000111111111100001111111100000000011", 
               "110000000000000000000000000000111111111110000000000000000000000000111111111000000000000001110000000000000011111111111111111111111000000000000001111111111111111111111110000000000000000000000000111111111111100000000000000000000000011111111110000000000000000000000000000111111111100001111111100000000011", 
               "110000111111100000001111110000000111110000000111111111111111110000000111111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110000000111111111111111110000000111111000000011111111111111111000000011111110000111111111111111111110000000011111100001111111100000000011", 
               "110000111111100000011111110000000111110000000111111111111111110000000111111000011111110000000000111111100000001111111111111111111000011111100000001111111111111111110000000111111111111111110000000111111000000011111111111111111000000011111110000111111111111111111110000000011111100001111111100000000011", 
               "110000111111100000011111110000000111110000000111111111111111110000000111111000011111110000000000111111100000001111111111111111111000011111100000001111111111111111110000000111111111111111110000000111111000000011111111111111111000000011111110000111111111111111111110000000011111100001111111100000000011", 
               "110000111111100000011111110000000111110000000111111111111111110000000111111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110000000111111111111111110000000111111000000011111111111111111000000011111110000111111111111111111110000000011111100001111111100000000011", 
               "110000111111100000011111110000000111110001111111100000000011111110000111111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110000111111100000000011111110000111111000000011111111111111111100000001111110000111111111111111111110000000011111100001111111100000000011", 
               "110000111111100000011111110000000111110001111111000000000001111110000000111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110001111111000000000001111111000000111000011111110000000000111111100000001110000000000011111100000000000000011111100001111111100000000011", 
               "110000111111100000011111110000000111110001111111000000000011111110000000111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110001111111000000000001111111000000111000011111110000000000111111100000001110000000000011111100000000000000011111100001111111100000000011", 
               "110000111111100000011111110000000111110001111111000000000011111110000000111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110001111111000000000001111111000000111000011111110000000000111111100000001110000000000011111100000000000000011111100001111111100000000011", 
               "110000111111100000011111110000000111110001111111000000000011111110000000111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110001111111000000000001111111000000111000011111110000000000111111100000001110000000000011111100000000000000011111100001111111100000000011", 
               "110000111111100000011111110000000111110001111111000000000011111110000000111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110001111111000000000001111111000000111000011111110000000000000000000000001111111111000011111100000000000000011111100001111111100000000011", 
               "110000111111100000011111110000000111110001111111000000000011111110000000111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110001111111000000000001111111000000111000011111110000000000000000000000001111111111000011111100000000000000011111100001111111100000000011", 
               "110000111111100000011111110000000111110001111111000000000001111110000000111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110001111111000000000001111111000000111000011111110000000000000000000000001111111111000011111100000000000000011111100001111111100000000011", 
               "110000111111100000011111110000000111110001111111000000000011111110000000111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110001111111000000000001111111000000111000011111110000000000000000000000001111111111000011111100000000000000011111100001111111100000000011", 
               "110000111111100000011111110000000111110001111111000000000011111110000000111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110001111111000000000001111111000000111000011111110000000000000000000000001111111111000011111100000000000000011111100001111100000000000011", 
               "110000000111111111111110000000000111110001111111000000000011111110000000111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110001111111000000000001111111000000111000000011111111111111111000000000001111111111000011111100000000111111111111100001111100000000000011", 
               "110000000111111111111110000000000111110001111111000000000011111110000000111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110001111111000000000001111111000000111000000011111111111111111000000000001111111111000011111100000001111111111111100001111100000000000011", 
               "110000000111111111111110000000000111110001111111000000000011111110000000111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110001111111000000000001111111000000111000000011111111111111111000000000001111111111000011111100000001111111111111100001111100000000000011", 
               "110000000111111111111110000000000111110001111111000000000011111110000000111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110001111111000000000001111111000000111000000011111111111111111000000000001111111111000011111100000000111111111111100001111100000000000011", 
               "110000000111111111111110000000000111110001111111000000000011111110000000111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110001111111000000000001111111000000111000000000011010000000111100100000001111111111000011111100000000111111111111100001111100000000000011", 
               "111111000000011111100000000000000111110001111111000000000011111110000000111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110001111111000000000001111111000000111000000000000000000000111111100000001111111111000011111100000001111111111111100001111100000000000011", 
               "111111000000011111100000000000000111110001111111000000000011111110000000111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110001111111000000000001111111000000111000000000000000000000111111100000001111111111000011111100000000111111111111100001111100000000000011", 
               "111111000000011111100000000000000111110001111111000000000011111110000000111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110001111111000000000001111111000000111000000000000000000000111111100000001111111111000011111100000000111111111111100001111100000000000011", 
               "111111000000011111100000000000000111110001111111000000000011111110000000111000011111110000000000111111100000011111111111111111111000011111100000001111111111111111110001111111000000000001111111000000111000000000000000000000111111100000001111111111000011111100000000111111111111100001111000000000000011", 
               "111111000000011111100000000000000111110001111111000000000011111110000000111000011111110000000000111111100000011111111111111111111000011111100000000000000000011111110001111111000000000001111111000000111000011111110000000000111111100000001111111111000011111100000000111111111111100001111100000000111111", 
               "111111111000011111100000000000111111110001111111000000000001111110000000111000011111110000000000111111100000011111111111111111111000011111100000000000000000011111110001111111000000000001111111000000111000011111110000000000111111100000001111111111000011111100000000111111111111100000000000000000111111", 
               "111111111000011111100000000000111111110001111111000000000011111110000000111000011111110000000000111111100000011111111111111111111000011111100000000000000000011111110001111111000000000001111111000000111000011111110000000000111111100000001111111111000011111100000000111111111111100000000000000000111111", 
               "111111111000011111100000000000111111110001111111000000000001111110000000111000011111110000000000111111100000011111111111111111111000011111100000000000000000011111110001111111000000000001111111000000111000011111110000000000111111100000001111111111000011111100000000111111111111100000000000000000111111", 
               "111111111000011111100000000000111111110000001111111111111111110000000000111000011111110000000000111111100000011111111111111111111000011111110000000000000000011111110000001111111111111111110000000000111000011111110000000000111111100000001111111111000011111100000000111111111111100000000000000000111111", 
               "111111111000011111100000001111111111110000000111111111111111110000000000111000000011111111111111111000000000011111111111111111111000011111111111111111111000000011110000000111111111111111110000000000111000000011111111111111111000000000001111111111000011111100000000111111111111100000000000000000111111", 
               "111111111000011111100000001111111111110000000111111111111111110000000000111000000011111111111111111000000000011111111111111111111000011111111111111111111000000011110000000111111111111111110000000000111000000011111111111111111000000000001111111111000011111100000000111111111111100001111100000000111111", 
               "111111111000011111100000001111111111110000000111111111111111110000000000111000000011111111111111111000000000011111111111111111111000011111111111111111111000000011110000000111111111111111110000000000111000000011111111111111111000000000001111111111000011111100000001111111111111100001111100000000111111", 
               "111111111000011111100000001111111111110000000111111111111111110000000000111000000011111111111111111000000000011111111111111111111000011111111111111111111000000011110000000111111111111111110000000000111000000011111111111111111000000000001111111111000011111100000000111111111111100001111100000000111111", 
               "111111111000011111100000001111111111110000000111111111111111100000000000111000000011111111111111111000000000011111111111111111111000011111111111111111111000000011110000000111111111111111110000000000111000000011111111111111111000000000001111111111000011111100000000111111111111100001111100000000111111", 
               "111111111000000000000000001111111111111110000000000000000000000000000000111111100000000000000000000000000000011111111111111111111000000000000000000000000000000011111110000000000000000000000000000000111111100000000000000000000000000000001111111111000000000000000000111111111111100001111100000000111111", 
               "111111111000000000000000001111111111111110000000000000000000000000000000111111100000000000000000000000000000011111111111111111111000000000000000000000000000000011111110000000000000000000000000000000111111100000000000000000000000000000001111111111000000000000000000111111111111100001111100000000111111", 
               "111111111000000000000000001111111111111110000000000000000000000000000000111111100000000000000000000000000000011111111111111111111000000000000000000000000000000011111110000000000000000000000000000000111111100000000000000000000000000000001111111111000000000000000000111111111111100001111000000000111111", 
               "111111111000000000000000001111111111111110000000000000000000000000000000111111100000000000000000000000000000011111111111111111111000000000000000000000000000000011111110000000000000000000000000000000111111100000000000000000000000000000001111111111000000000000000000111111111111100000000000000000111111", 
               "111111111000000000000000001111111111111111110000000000000000000000000111111111100000000000000000000000000000011111111111111111111111000000000000000000000000000011111111111000000000000000000000000111111111111100000000000000000000000001111111111111111100000000000000111111111111100000000000000000111111", 
               "111111111111100000000000001111111111111111110000000000000000000000000111111111111100000000000000000000000011111111111111111111111111100000000000000000000000000011111111111000000000000000000000000111111111111100000000000000000000000011111111111111111100000000000000111111111111100000000000000000111111", 
               "111111111111100000000000001111111111111111111000000000000000000000000111111111111100000000000000000000000011111111111111111111111111100000000000000000000000000011111111111000000000000000000000000111111111111100000000000000000000000011111111111111111100000000000000111111111111100000000000000000111111", 
               "111111111111100000000000001111111111111111110000000000000000000000000111111111111100000000000000000000000011111111111111111111111111000000000000000000000000000011111111111000000000000000000000000111111111111100000000000000000000000011111111111111111100000000000000111111111111100000000000000000111111", 
               "111111111111100000000000001111111111111111111000000000000000000000000111111111111100000000000000000000000011111111111111111111111111100000000000000000000000000011111111111000000000000000000000000111111111111100000000000000000000000011111111111111111100000000000000111111111111111110000000000000111111", 
               "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111", 
               "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111", 
               "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111", 
               "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111", 
               "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111", 
               "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
               "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");
            
 GS_message <= ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1110000000000000001111110000000000000000111111000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1110000000000000000111110000000000000000111111000000000000000001111111000000000000001111111100000000000000111111111111111111111111110000000000001111111100000000000000001111111111111111111111111111111111111111111111111111111111111111111100000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1110000000000000000111110000000000000000111111000000000000000000111111000000000000001111111100000000000000111111111111111111111111100000000000000111111000000000000000000111000000001100000000111000000000000000011110000000000000000001111100000000000000011111111111111111111111100000000000000001111111111111111111111111111100000000000000011100000000000000001111110000000000000111111110000001110000000111",
                "1110011111111111000011110001111111111000011111001111111111111000011110000000000000001111111000000000000000011111111111111111111111100000000000000111111000000000000000000111000000001100000000111000000000000000011110000000000000000001111100000000000000001111111111111111111111100000000000000001111110000000011000000011111000000000000000011100000000000000001111100000000000000111111100000000110000000111",
                "1110011111111111100001110011111111111100001111001111111111111100011100001111111111000011110000111111111000011111111111111111111111000011111111000011111000111111111111000111000000001100000000111000000000000000011110000000000000000001111100111111111110000111111111111111111111100000000000000001111110000000011000000001111000000000000000011100000000000000001111100000000000000011111100000000110000000011",
                "1110011111111111100001110011111111111100001111001111111111111000011100001111111111000011110000111111111100001111111111111111111110000111111111100001111001111111111111100011001111000000111100001001111111111110000110001111111111111000111000111111111110000111111111111111111111100111111111110000011110000000010000000001111000111111111100001100111111111111000110000111111111100001111100011000000011100001",
                "1110011110000001111000110011110000001111000111001111000000000000011100011110000111100001110001110000011110000111111111111111111110000111111111100001111001111111111111100011001111000000111100001001111111111110000110001111111111111000011100111111111111000011111111111111111111100111111111111000011110011110000001111000111001111111111110000100111111111111000010000111111111100001111100111100000011110001",
                "1110011110000001111000110011110000001111000011001111000000000000011100111100000011110001110011110000001111000111111111111111111110001111000001111000111001111000000000000011001111100000111100001000111111111100000110001111111111111000011100111100000111100001111111111111111111100111111111111000011110011110000001111000111001111111111110000100011111111110000010001111000011110000111100111100000011110001",
                "1110011110000001111000110011110000001111000011001111000000000000011100111100000011110001110011110000001111000111111111111111111110001110000001111000011001111000000000000011001111110000111100001000000111100000000110001111000000000000011100111100000011100001111111111111111111100111100000011110001110011110000001111000111000000111100000000100000011110000000010001110000001111000011100111110000011110001",
                "1110011110000001111000110011110000001111000011001111000000000000011100111100000000000001110011110000000000000111111111111111111110011110000000111000011001111000000000000011001111111000111100001100000111100000000110001110000000000000011100111100000011110001111111111111111111100111100000011110000110011110000001111000111000000111100000000100000011110000000010011110000001111000011100111111000011110001",
                "1110011110000001111000110011111000001111000011001111000000000000011100111100000000000001110011110000000000000111111111111111111110001110000000000000011001111000000000000011001111111100111100001111100111100000000110001110000000000000011100111100000011100001111111111111111111100111100000011110000110011110000001111000111100000111100000000111100011110000000010011110000001111000011100111111000011110001",
                "1110011110000001111000110011111111111100000011001111111111100000111100011100000000000001110011110000000000000111111111111111111110011110000000000000011001111000000000000011001111111100111100001111100111100000000110001111000000000000111100111100000111100001111111111111111111100111100000011110001110011110000001111000111111100111100000000111110011110000000010011110000001111000011100111111100011110001",
                "1110011110000001111000110011111111111100000011001111111111100001111100001111111111000001110000111111111000000111111111111111111110001110000000000000011001111111111100000111001111111100111100001111100111100000000110001111000000000000111100111111111110000001111111111111111111100111100000111100001110011110000001111000111111100111100000000111110011110000000110011110000001111000011100111111100011110001",
                "1110011111000011110000110011111111111110000011001111111111100001111100001111111111000001110000111111111100000111111111111111111110011110000000000000011001111111111110000111001111001111111100001111100111100001111110001111111111100001111100111111111110000001111111111111111111100111111111111000001110011110000001111000111111100111100000101111110011110000111110011110000001111000011100111101110111110001",
                "1110011111111111100000110011110000001111000011001111000000000001111100000111111111000001110000011111011100000111111111111111111110011110000000000000011001111111111100000111001111001111111100001111100111100001111110001111111111100001111100111111111110000001111111111111111111100111111111111000001110011110000001111000111111100111100001111111110011110000111110011110000001111000011100111100111111110001",
                "1110011111111111100000110011110000001111000011001111000000000001111100000000000011110001110000000000001111000111111111111111111110001110000000000001111001111000000000000111001111000011111100001111100111100001111110001111000000000001111100111100000111100001111111111111111111100111100000111100001110011110000001111000111111100111100001111111110011110000111110001110000001111000011100111100111111110001",
                "1110011111111111000000110011110000001111000011001111000000000001111100000000000011110001110000000000001111000111111111111111111110001110000000000001111001111000000000000111001111000011111100001111100111100001111110001111000000000001111100111100000011110001111111111111111111100111100000011110001110011110000001111000111111100111100001111111110011110000111110011110000001111000011100111100011111110001",
                "1110011110000000000000110011110000001111000011001111000000000001111100011100000011110001110011100000001111000111111111111111111110001110000000000001111001111000000000000111001111000011111100001111100111100001111110001111000000000001111100111100000011100001111111111111111111100111100000011110001110011110000001111000111111100111100001111111110011110000111110011110000001111000011100111100001111110001",
                "1110011110000000000000110011110000001111000011001111000000000000111100111100000011110001110011110000001111000111111111111111111110001110000001111000011001111000000000000111001111000000111100001111100111100001111110001110000000000001111100111100000011100001111111111111111111100111100000011110000110011110000001111000111111100111100001111111110011110000111110011110000001111000011100111100001111110001",
                "1110011110000000000001110011110000001111000011001111111111111000011100011110000011100001110001111000011110000111111111111111111110001110000001111000011001111000000000000111001111000000111100001111100111100001111110001110000000000001111100111100000011100001111111111111111111100111100000011110001110011110000001111000111111100111100001111111110011110000111110001110000001111000011100111100000111110001",
                "1110011110000000000001110011110000001111000011001111111111111100011100001111111111000001110000111111111100000111111111111111111110001111000001111000011001111100111001000111001111000000111100001111100111100001111110001111000000000001111100111100000011100001111111111111111111100111100000011100000110011110000001111000111111100111100001111111110011110000111110001111000001111000011100111100000011110001",
                "1110011110000000000011110001110000001111000011001111111111111100011100001111111111000001110000111111111100000111111111111111111110000111111111100000011001111111111111100011001111000000111100001111100111100001111110001111111111111000111000111100000111100001111111111111111111100111111111111000000110011110000011110000111111100111100001111111110011110000111110000111111111100000011100111100000011110001",
                "1110000000000111111111110000000000000000000011000000000000000000011110001111111110000001110000111111111000000111111111111111111110000111111111100000011001111111111111100011001111000000111100001111100111100001111110001111111111111000011000111000000011100001111111111111111111100111111111111000001110000111111111100000111111100111100001111111110011110000111110000111111111100000011100111100000011110001",
                "1110000000000111111111110000000000000000000011000000000000000000011111000000000000000001111100000000000000000111111111111111111111000011111111000000011000111111111111000011000111000000011100001111100011100001111110001111111111111000011100000000000000000001111111111111111111100111111111110000000110000111111111100000111111100111100001111111110011100000111111000011111111100000011100111100000011110001",
                "1110000000000111111111111000000000000000000011000000000000000000011111000000000000000001111100000000000000000111111111111111111111100000000000000000011000000000000000000011000000000000000000001111100000000001111110000000000000000000011100000000000000000001111111111111111111100000000000000000000110000111111111000000111111100000000001111111110000000000111111100000000000000000011100011000000010000001",
                "1111100000000111111111111100000000110000000011110000000000000000011111100000000000000011111110000000000000001111111111111111111111110000000000000000011000000000000000000011000000000000000000001111100000000001111110000000000000000000011100000000000000000001111111111111111111100000000000000000001111100000000000000000111111100000000001111111110000000000111111110000000000000000011100000000000000000001",
                "1111100000000111111111111100000000110000000011110000000000000000011111110000000000000011111111000000000000001111111111111111111111111000000000000000111110000000000000000011100000000000000000001111110000000001111111000000000000000000011110000000001000000001111111111111111111110000000000000000001111100000000000000000111111100000000001111111110000000000111111110000000000000000111100000000000000000001",
                "1111110010001111111111111110001001111000000111110000000000000000011111110000000000000011111111000000000000001111111111111111111111111000000000000001111110000000000000000011110000000011000000001111111000000001111111100000000000000000011111000000011100000001111111111111111111111000000000000000011111110000000000000000111111111000000001111111111100000000111111111000000000000001111110000000001000000001",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000001111110000000000000000011111000000011000000001111111000000001111111110000000000000000111111000000011100000001111111111111111111111000000000000000111111111000000000000001111111111000000001111111111100000000111111111000000000000001111111000000001100000001",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000011111111111100000011111111111111111111111111111111111111111111111111000000011100000001",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",         
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111100000000000001111111111111111111111110111111111111111110000000000000001111111000000000000011111110000000000000000111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011111100000000000000111111111111111111111100000000000000111110000000000000001111111000000000000001111110000000000000000111111000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000011111100000000000000111111111111111111111100000000000000111110000000000000000111110000000000000001111110000000000001000011111001111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000111111111100001110000111111111000011111111111111111111000000000000000011110011111111111000011100001111111110000111110011111111111100001111001111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111110000110000111111111000011111111111111111110000111111111100001100011111111111000011100001111111111000011110011111111111100001111001111111111100001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001111111111100000110001111111111100001111111111111111110000111111111100001110011111111111000011100011110000111100011110011111000001110000111000000111000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111100000000110011110000001110000111111111111111110001111000001111000110000001111000000011100111100000011100001110011110000001111000011000000111000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111100000000110011110000001111000111111111111111110011110000001111000110000001110000000011100111100000011110001110011110000001111000011110000111000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000111100000000110011110000001111000111111111111111110011110000001111000110000001110000000011100111100000011110001110011110000001111000011111100111000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111100000000110011110000001111000111111111111111110011110000000000000111110001110000000011100111100000011110001110011110000001111000011111100111000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111100000000110011110000001111000111111111111111110011110000000000000111111001110000000011100111100000011110001110011111000011110000011111100111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111100001101110011110000001111000111111111111111110001110000000000000111111001110000011111100111100000011110001110011111111111100000011111100111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111100001111110011110000001111000111111111111111110000111111111100000111111001110000111111100111100000011110001110011111111111100000011111100111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111100001111110011110000001111000111111111111111110000111111111100000111111001110000111111100111111111111110001110011111000001110000011111100111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111100001111110011110000001111000111111111111111110000011111111110000111111001110000111111100111111111111110001110011110000001111000011111100111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111100001111110011110000001111000111111111111111110000000000001111000111111001110000111111100111111111111110001110011110000001111000011111100111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111100001111110011110000001111000111111111111111110000000000001111000111111001110000111111100111100000111110001110011110000001111000011111100111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111100001111110011110000001111000111111111111111110001110000001111000111110001110000111111100111100000011110001110011110000001111000011111100111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111100001111110011110000001110000111111111111111110011110000001111000111111001110000111111100111100000011110001110011110000001111000011111100111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111100001111110001111111111100000111111111111111110001111000001110000111111001110000111111100111100000011110001110011110000001111000011111100111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111100001111110000111111111000000111111111111111110000111111111100000111110001110000111111100111100000011100001110011110000001111000011111100111000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100111100001111110000111111111000000111111111111111110000111111111100000111110001110000111111100111000000011100001110001110000000110000011111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111111000000000000000000111111111111111111000011111111000000111111000000000111111100000000000000000001110000000000000000000011111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111111100000000000000000111111111111111111100000000000000000111111000000000111111100000000000000000001110000000000000000000011111100000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111111100000000000000000111111111111111111100000000000000000111111000000000111111110000000001000000001111100000000110000000011111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000001111111110000000000000001111111111111111111111000000000000001111111100000000111111111000000011100000001111100000000110000000011111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000001111111111000000000000011111111111111111111111000000000000001111111110000000111111111000000011100000001111110000000110000000111111111000110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011111111111000000000000011111111111111111111111000000000000001111111110000000111111111110111111100111001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");
                                                                                                                                                                                                                                                                                                                                                                                                                                 
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
   
IngameLogoTop <=("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000011111111111111111111111111111111000000000010011111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000011111111111111111111111111000000000000000000000000011111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000111111111111111111111110000000000000000000000000000000001111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000001111111111111111111110000000000000000000000000000000000000001111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000111111111111111111110000000000000000000000000000000000000000000011111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000001111111111111111110000000000000000000000000000000000000000000000000011111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111111111111111100000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000111111111111111111111111111",
                 "11111111111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111",
                 "11111111111111111111111111111111111111111100000000000000000000000000000001111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
                 "11111111111111111111111111111111111111000000000000000000000000000000000000001111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
                 "11111111111111111111111111111111111100000000000000000000000000000000000000000001111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
                 "11111111111111111111111111111111100000000000000000000000000000000000000000000000011111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
                 "11111111111111111111111111111110000000000000000000000000000000000000000000000000000011111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111",
                 "11111111111111111111111111111000000000000000000000000000000000000000000000000000000000111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111",
                 "11111111111111111111111111100000000000000000000000000000000000000000000000000000000000011111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111",
                 "11111111111111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111",
                 "11111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111",
                 "11111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000011111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111",
                 "11111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000001111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111",
                 "11111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111",
                 "11111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111",
                 "11111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111",
                 "11111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111",
                 "11111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111",
                 "11111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111",
                 "11111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111",
                 "11111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111",
                 "11111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111",
                 "11111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
                 "11111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
                 "11111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
                 "11111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
                 "11111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
                 "11111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
                 "11111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
                 "11111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
                 "11111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
                 "11111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
                 "11111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111",
                 "11111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111",
                 "11111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111",
                 "11111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111",
                 "11111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111",
                 "11111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111",
                 "11111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111",
                 "11111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111",
                 "11111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111",
                 "11111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111",
                 "11110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111",
                 "11110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111",
                 "11110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111",
                 "11110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111",
                 "11110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111",
                 "11110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111",
                 "11110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111",
                 "11110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
                 "11110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
                 "11110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
                 "11110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111",
                 "11110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
                 "11110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
                 "11111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
                 "11111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111",
                 "11111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
                 "11111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111",
                 "11111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111",
                 "11111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111",
                 "11111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111",
                 "11111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111",
                 "11111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111",
                 "11111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111",
                 "11111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111",
                 "11111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111",
                 "11111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110000000000000000000000000000000000000000000000000000000000000000000000000111111111111",
                 "11111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000000000000000001111111111111",
                 "11111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000001111111110000000000000000000000000000000000000000000000000000000000000000011111111111111",
                 "11111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111100000000001111111111110000000000000000000000000000000000000000000000000000000000000011111111111111",
                 "11111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111100000000011111111111111110000000000000000000000000000000000000000000000000000000000111111111111111",
                 "11111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111000000000011111111111111111110000000000000000000000000000000000000000000000000000001111111111111111",
                 "11111111111000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111000000000111111111111111111111110000000000000000000000000000000000000000000000000011111111111111111",
                 "11111111111100000000000000000000000000000000000000000000000000000000000000000000000000011111111111110000000000111111111111111111111111110000000000000000000000000000000000000000000000111111111111111111",
                 "11111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111111100000000001111111111111111111111111111110000000000000000000000000000000000000000001111111111111111111",
                 "11111111111110000000000000000000000000000000000000000000000000000000000000000000001111111111111111100000000000111111111111111111111111111111110000000000000000000000000000000000000011111111111111111111",
                 "11111111111111000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000001111111111111111111111111111111110000000000000000000000000000000000111111111111111111111",
                 "11111111111111100000000000000000000000000000000000000000000000000000000000000111111111111111111110000000000000000011111111111111111111111111111111110000000000000000000000000000001111111111111111111111",
                 "11111111111111100000000000000000000000000000000000000000000000000000000000111111111111111111111100000000000000000001111111111111111111111111111111111110000000000000000000000000011111111111111111111111",
                 "11111111111111110000000000000000000000000000000000000000000000000000000111111111111111111111111000000000000000000000111111111111111111111111111111111111110000000000000000000001111111111111111111111111",
                 "11111111111111111000000000000000000000000000000000000000000000000000011111111111111111111111110000000000000000000000011111111111111111111111111111111111111100000000000000000011111111111111111111111111",
                 "11111111111111111100000000000000000000000000000000000000000000000011111111111111111111111111100000000000100000000000011111111111111111111111111111111111111100000000000000000111111111111111111111111111",
                 "11111111111111111110000000000000000000000000000000000000000000011111111111111111111111111111000000000001111000000000111111111111111111111111111111111111100000000000000000011111111111111111111111111111",
                 "11111111111111111111000000000000000000000000000000000000000011111111111111111111111111111100000000000011111000000000111111111111111111111111111111110000000000000000000000111111111111111111111111111111",
                 "11111111111111111111100000000000000000000000000000000000001111111111111111111111111111111000000000000111111000000000111111111111000000000000000000000000000000000000000011111111111111111111111111111111",
                 "11111111111111111111110000000000000000000000000000000001111111111111111111111111111111100000000000001111110000000001111111111110000000000000000000000000000000000000001111111111111111111111111111111111",
                 "11111111111111111111111100000000000000000000000000001111111111111111111111111111111111000000000000011111110000000001111111111110000000000000000000000000000000000000111111111111111111111111111111111111",
                 "11111111111111111111111110000000000000000000000000111111111111111111111111111111111110000000000000111111100000000011111111111100000000000000000000000000000000000111111111111111111111111111111111111111",
                 "11111111111111111111111111000000000000000000000111111111111111111111111111111111111110000000000001111111100000000011111111111100000000000000000000000000000000111111111111111111111111111111111111111111",
                 "11111111111111111111111111110000000000000000001111111111111111111111111111111111111110000000000111111111000000000111111111111000000000000000000000000000000111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111000000000000000000111111111111111111111111111111111111111000000000111111111000000000111111111111000000000000000000000000001111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111110000000000000000000001111111111111111111111111111111111000000000111111110000000000111111111111000000000000000000011111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111000000000000000000000000000111111000000000111111111111100000000011111110000000001111111111110000000001111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111110000000000000000000000000000000000000000011111111111100000000011111100000000001111111111110000000001111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111100000000000000000000000000000000000000011111111111110000000001111100000000011111111111100000000011111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111100000000000000000000000000000000000001111111111110000000001111100000000011111111111100000000011111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111100000000000000000000000000000000001111111111110000000000111000000000111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111100000000000000000000000000000000111111111111000000000111000000000111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111110000000000000000000000000000111111111111100000000010000000001111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111100000000000000000000000011111111111100000000000000000001111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111100000000011111111111110000000000000000011111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111110000000001111111111110000000000000000011111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111110000000001111111111111000000000000000111111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111000000000000000111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111100000000000000111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111100000000000001111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111110000000000001111111111110000000001111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111110000000001111111111110000000000011111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111110000000001111111111110000000000001111111111100000000011111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111000000000000001111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111000000000000000001111000000000111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111100000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111100000000011111111111100000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111100000000001111111111110000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111110000000001111111111110000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111110000000000111111111110000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111110000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111100000000011111000000000000000011000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111100000000001000000000000000000111111000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000111111111000011111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111110000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"); 

IngameLogoBottom <=( "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110001111111110000000000011111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000011111111110000000000000011111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000111111111100000000000000000111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111100000000000000000000011111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000001111111111000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000001111111111000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000001111111111000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000111111111111100000000000000000000000000000000111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000001111111111111111000000000000000000000000000000000111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000011111111111111111100000000000000000000000000000000000011111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000111111111111111111111000000000000000000000000000000000000011111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000001111111111111111111111100000000000000000000000000000000000000111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000011111111111111111111111110000000000000000000000000000000000000001111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000111111111111111111111111110000000000000000000000000000000000000001111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111000000000000000000000000000001111111111111111111111111100000000000000000000000000000000000000011111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111100000000000000000000000000000000111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111000000000000000000000000000000001111111111111111111111111111000000000000001111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111000000000000000000000000000000000011111111111111111111111111111000000000000011111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111110000000000000000000000000000000000011111111111111111111111111110000000000000111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111110000000000000000000000000000000000001111111111111111111111111111110000000000000111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111100000000000000000000000000000000000000011111111111111111111111111111100000000000001111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111000000000000000000000000000000000000000011111111111111111111111111111100000000000001111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111000000000000000000000000000000000000000001111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111100000000000000000000000000000000000001111111111111111111111111111000000000000011111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111110000000000111100000000000000111111111111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111000000000000011111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111000000000000111111111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111000000000000111111111111111111111000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000011111111111110000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000111111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                     "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");                  
                     
                     
                 
    PongNameLabel <= ("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000011111111111111110000000000000000000000111110000000000000000000000011111111111111100000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000011111111111111110000000000000000000000111110000000000000000000000011111111111111100000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000011111111111111110000000000000000000000111110000000000000000000000011111111111111100000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000011111111111111110000000000000000000000111110000000000000000000000011111111111111100000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000011111111111111110000000000000000000000111110000000000000000000000011111111111111100000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000011111111111111111111100000000000000000000000000000000000000011111111111111110000000000000000000000111110000000000000000000000011111111111111100000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000001111111111111111111100000000000000000000000000000000000000011111111111111110000000000000000000000111110000000000000000000000011111111111111100000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111111111111111111111111100000000000011111111100000000000111111111111111111111111111100000000000111111111110000001111111111100000000000000001111111111100000000000111100000000000111111111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111111111111111111111111100000000000011111111100000000000111111111111111111111111111100000000000111111111110000001111111111100000000000000001111111111100000000000111100000000000111111111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111111111111111111111111100000000000011111111100000000000111111111111111111111111111100000000000111111111110000001111111111100000000000000001111111111100000000000111100000000000111111111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111111111111111111111111100000000000011111111100000000000111111111111111111111111111100000000000111111111110000001111111111100000000000000001111111111100000000000111100000000000111111111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111111111111111111111111100000000000011111111100000000000111111111111111111111111111100000000000111111111110000001111111111100000000000000001111111111100000000000111100000000000111111111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111111111111111111111111100000000000011111111100000000000111111111111111111111111111100000000000111111111110000001111111111100000000000000001111111111100000000000111100000000000111111111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111111111000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111111111000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111111111000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111111111000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111111111000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111111111111110000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111111111111110000001111111111100000000000111100000011111111111000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111111111111110000001111111111100000000000111100000011111111111000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111111111111110000001111111111100000000000111100000011111111111000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111111111111110000001111111111100000000000111100000011111111111000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111111111111110000001111111111100000000000111100000011111111111000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111111111111110000001111111111100000000000111100000011111111111000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111100000111111111111111111111100000000000111100000011111111111000000000001111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111100000111111111111111111111100000000000111100000011111111111000000000001111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111100000111111111111111111111100000000000111100000011111111111000000000001111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111100000111111111111111111111100000000000111100000011111111111000000000001111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111100000111111111111111111111100000000000111100000011111111111000000000001111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111100000111111111111111111111100000000000111100000011111111111000000000001111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111111111111111111111111100000000000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111100000000001111111111111111100000000000111100000011111111111000000000000000001111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111111111111111111111111100000000000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111100000000001111111111111111100000000000111100000011111111111000000000000000001111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111111111111111111111111100000000000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111100000000001111111111111111100000000000111100000011111111111000000000000000001111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111111111111111111111111100000000000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111100000000001111111111111111100000000000111100000011111111111000000000000000001111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111111111111111111111111100000000000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111100000000001111111111111111100000000000111100000011111111111000000000000000001111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111111111111111111111111100000000000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111100000000001111111111111111100000000000111100000011111111111000000000000000001111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000000000000000000000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111100000000000100001111111111100000000000111100000011111111111000000000000000001111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000000000000000000000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000000000000000000000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000000000000000000000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000000000000000000000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111100000000000000001111111111100000000000111100000011111111111000000000000000001111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000000000000000000000000000111100000011111111111000000000000000001111111111100000000001111110000001111111111100000000000000001111111111100000000000111100000011111111111100000000000000001111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000000000000000000000011111111100000000000111111111111111111111111111100000000000000001111110000001111111111100000000000000001111111111100000000000111100000000000111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000000000000000000000011111111100000000000111111111111111111111111111100000000000000001111110000001111111111100000000000000001111111111100000000000111100000000000111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000000000000000000000011111111100000000000111111111111111111111111111100000000000000001111110000001111111111100000000000000001111111111100000000000111100000000000111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000000000000000000000011111111100000000000111111111111111111111111111100000000000000001111110000001111111111100000000000000001111111111100000000000111100000000000111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000000000000000000000011111111100000000000111111111111111111111111111100000000000000001111110000001111111111100000000000000001111111111100000000000111100000000000111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111100000000000000000000000000000000011111111100000000000111111111111111111111111111100000000000000001111110000001111111111100000000000000001111111111100000000000111100000000000111111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000101110000000000000000111111111100000000000011111111111111111111111111100000000000000001111110000000000000000000000000000000000000000000000000000000111100000000000011111111111111111111111111111111100000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000001111111111111111111111111111111111111100000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000111111111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000001111111111111111111111111111111111111110000000000000000000000000000000000000000000000001111110000000000000000000000000000000000000000000000000000000111111111110000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000000000111111111111111100000000000000000000001111110000000000000000000000111111111111111000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000000000111111111111111100000000000000000000001111110000000000000000000000111111111111111000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000000000111111111111111100000000000000000000001111110000000000000000000000111111111111111000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000000000111111111111111100000000000000000000001111110000000000000000000000111111111111111000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000000000111111111111111100000000000000000000001111110000000000000000000000111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000001111111111111111111111111111111111111111111000000000000000000000000000000000000000111111111111111110000000000000000000001111110000000000000000000000111111111111111000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111",
                  "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");


    ponglogo <=("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111000000000000000111111111111111111111111111101111011111111111111110000000001111111111100001111111111100011111111111000000000111111111111111111",
                "1111111111111111111000000000000000111111111111111111111111100000000000011111111111100000000000111111111100001111111111000011111111110000000000011111111111111111",
                "1111111111111111111000000000000000111111111111111111111111000000000000001111111111000000000000011111111100000111111111000011111111100000000000001111111111111111",
                "1111111111111111111000000000000000011111111111111111111111000000000000000111111111000000000000001111111000000111111111000011111111000000000000000111111111111111",
                "1111111111111111000000000000000000000011111111111111111111000000000000000111111110000000000000001111111000000111111111000011111111000000000000000111111111111111",
                "1111111111111111000000000000000000000011111111111111111111000000000000000011111100000000000000000111111000000011111111000011111110000000000000000011111111111111",
                "1111111111111111000000000000000000000011111111111111111111000000000000000011111100000011111000000111111000000011111111000011111110000001111100000011111111111111",
                "1111111111111111000000000000000000000011111111111111111111000011111100000011111100000111111100000011111000000011111111000011111100000011111110000001111111111111",
                "1111111111111111000000000000000000000011111111111111111111000011111110000011111000000111111100000011111000000001111111000011111100000111111110000001111111111111",
                "1111111111111111000000000000000000000011111111111111111111000011111111000001111000001111111110000011111000000001111111000011111100000111111111000001111111111111",
                "1111111111111110000000000000000000000011111111111111111111000011111111000001111000001111111110000001111000000001111111000011111000001111111111000001111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111000001110000011111111111000001111000000000111111000011111000001111111111100001111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111000001110000011111111111000001111000000000111111000011111000001111111111100001111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111000001110000011111111111000001111000000000011111000011111000001111111111100011111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111000001110000011111111111000001111000000000011111000011111000011111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111000001110000011111111111100001111000000000011111000011110000011111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111000001110000111111111111100001111000001000001111000011110000011111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111110000011110000111111111111100000111000001000001111000011110000011111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111100000011110000111111111111100000111000001000001111000011110000011111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111000000000000000011110000111111111111100000111000001100000111000011110000011111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111000000000000000011110000111111111111100000111000001100000111000011110000011111110000000011111111111111",
                "1111111111110000000000000000000000000000001111111111111111000000000000000111110000111111111111100000111000001100000111000011110000011111110000000001111111111111",
                "1111111111110000000000000000000000000000001111111111111111000000000000000111110000111111111111100000111000001110000011000011110000011111100000000001111111111111",
                "1111111111110000000000000000000000000000001111111111111111000000000000001111110000111111111111100000111000001110000011000011110000011111100000000000111111111111",
                "1111111111110000000000000000000000000000001111111111111111000000000000011111110000111111111111100000111000001110000011000011110000011111100000000000111111111111",
                "1111111111110000000000000000000000000000001111111111111111000000000001111111110000111111111111100001111000001111000001000011110000011111110000000000111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111111111110000011111111111100001111000001111000001000011110000011111111111100000111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111111111110000011111111111000001111000001111100001000011111000011111111111100000111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111111111110000011111111111000001111000001111100000000011111000001111111111100000111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111111111110000011111111111000001111000001111100000000011111000001111111111100000111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111111111110000011111111111000001111000001111110000000011111000001111111111100000111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111111111111000001111111110000001111000001111110000000011111000001111111111100000111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111111111111000001111111110000011111000001111110000000011111100000111111111100000111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111111111111000000111111110000011111000001111111000000011111100000111111111100000111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111111111111100000111111100000011111000001111111000000011111100000011111111000000111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111111111111100000011111000000111111000001111111000000011111110000001111110000001111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111111111111100000000000000000111111000001111111100000011111110000000000000000001111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111111111111110000000000000001111111000001111111100000011111111000000000000000001111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111111111111110000000000000001111111000001111111100000011111111000000000000000011111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111111111111111000000000000011111111000001111111110000011111111100000000000000111111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111111111111111100000000000111111111100011111111110000011111111110000000000001111111111111111",
                "1111111111110000000000000000000000000000001111111111111111000011111111111111111111110000000001111111111100011111111111000111111111111000000000111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111100111111111111111111111111100000111111111111110111111111111100111111111111110000011111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111110000000000000001111000000000000000111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111110000000000000001111000000000000000111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111110000000000000001111000000000000000111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111110000000000000001111000000000000000111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111110000000000000001111000000000000000111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111110000000000000001111000000000000000111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111110000000000000001111000000000000000111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000011111111111111110011111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000011111111111111100011111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000011111111111111100011111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000011111111111111100011111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000011111111111111100011111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000011111111111111100011111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000011111111111111110011111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111100000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000000000000000000000001111111110000000001111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000011111111111111100011111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000011111111111111100011111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000011111111111111100011111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000011111111111111100011111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000011111111111111100011111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000011111111111111100011111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000011111111111111110011111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111110000000000000001111000000000000000111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111110000000000000001111000000000000000111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111110000000000000001111000000000000000111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111110000000000000001111000000000000000111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111110000000000000001111000000000000000111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111110000000000000001111000000000000000111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111110000000000000001111000000000000000111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111110000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111011000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111100000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");
                
                
                
 ArrowLogo_Name <=
("1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111100000000000011100000000000011100000010000001111000001100000011000000011111000000000011111111",
 "1111111000000000001100000000000001111000000000000111100000010000000100000000000001100000000000011100000010000000110000000100000011000000011111000000000001111111",
 "1111111000000000001100000000000001111000000000000111100000010000000100000000000011100000000000011100000010000001110000000100000011000000011111000000000011111111",
 "1111111000000000001100000000000001111000000000000111100000010000000100000000000000100000000000001100000000000000010000000000000001000000001100000000000000111111",
 "1111100001111110000100011111111000111001111111100011100110000011000000111000111000100111111110000100110000011100010011100000110001001110001100011111110000111111",
 "1111100001111110000100011111111000111001111111100011100110000011100000111000110000100111111110000100110000011100010001100000110001000110001100001111110000111111",
 "1111100011000010000100011100011000011001110001100001100110000011100000111000110000100000110000000100110000011100010001100001110001000110001100011000011000011111",
 "1111100111000001100100011000001100011001100000110000100110000011100000111000110000100000110000000100110000011100010001110011110001000110001100110000001100011111",
 "1111100111000001100100011000001100001001100000110000100110000011100000111000110000100000110000000100110000011100010001110011110001000110001100111000001100011111",
 "1111100111000001100100011000001100011001100000110000100110000011100000111000110000111100110000000100110000011100010001111111110001000110001100111000001100011111",
 "1111100111000001100100011000001100011001100000110000100110000011100000111000110000111100110000000100110000011100010001111111110001000110001100111000001100011111",
 "1111100111000001100100011000001100011001100000110000100110000011100000011000110000111100110000000100110000011100010001101101110001000110001100111000001100011111",
 "1111100111000001100100011000011000011001110001100000100111000011100000001111100000111100110000111100111111111100010001100100110001000110001100111000001100011111",
 "1111100111000001100100011111111000011001111111100000100111111111100000001111100000111100110000111100111111111100010001100100110001000110001100111000001100011111",
 "1111100111000001100100011100011000011001110001100000100111000011100010000111000000111100110000111100110000011100010001100000110001000110001100111000011100011111",
 "1111100111111111100100011000001100011001100000110000100110000011100011000110000000111100110000111100110000011100010001100000110001000110001100111111111100011111",
 "1111100111111111100100011000001100011001100000110000100110000011100011000110000000111100110000111100110000011100010001100000110001000110001100111111111100011111",
 "1111100111000011100100011000001100011001100000110000100110000011100011000110000000111100110000111100110000011100010001100000110001000110001100111000011100011111",
 "1111100111000001100100011000001100011001100000110000100110000011100011100110000001111100110000111100110000011100010001100000110001000110001100110000001100011111",
 "1111100111000001100100011000001100011001100000110000100110000011100011100110000001111100110000111100110000011100010001100000110001000110001100111000001100011111",
 "1111100111000001100100011000001100011001100000110000100110000011100011100110000111111100110000111100110000011100010001100000110001000110001100111000001100011111",
 "1111100111000001100100011000001100011001100000110000100110000011100011100110000111111100110000111100110000011100010001100000110001000110001100111000001100011111",
 "1111100111000011100100011000001100011001100000111000100110000011100011100110000111111100110000111100110000011000010001100000110001000110001100110000001100011111",
 "1111100000000000000100000000000000011000000000000000100000000000000011100000000111111100000000111100000000000000010000000000000001000000001100000000000000011111",
 "1111100000000000000100000000000000011000000000000000100000000000000011100000000111111100000000111100000000000000010000000000000001000000001100000000000000011111",
 "1111100000000000000100000000000000011000000000000000100000000000000011100000000111111100000000111100000000000000011000000000000001000000001100000000000000011111",
 "1111110000000100000111000000100000001100000000000000110000000100000011111000000111111110000000111110000001100000011100000010000000110000001111000000100000011111",
 "1111111000000100000111000000110000001100000011000000110000001100000011111000000111111110000000111110000001100000011100000010000000110000001111000000100000011111",
 "1111111000000100000111000000100000001100000011000000110000001100000011111000000111111110000001111111000001100000011100000010000001110000001111000000100000011111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");
               
                
    
  Arrowlogo <=( "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111001111111110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111110000111111110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111100000011111110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111000000001111110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111110000000000111110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111100000000000011110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111100000000000011110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111110000000100111110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111010000111111110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111110000111111110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111110000111111110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111001111111110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111111111111110001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111110000000000000000000000011111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111",
                "1111111111111111111111100000000000000000000000001111111111111111111111111111111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
                "1111111111111111111111000000000000000000000000000111111111111111111111111111111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
                "1111111111111111111111000111111111111111111110000111111111111111111111111111111111111111111111111111111110001111111111111111111100011111111111111111111111111111",
                "1111111111111111111111000111111111111111111110000111111111111111111111111111111111111111111111111111111110001111111111111111111100011111111111111111111111111111",
                "1111111111111111111111000111111111111111111110000111111111111111111111111111111111111111111111111111111110001111111111111111111100011111111111111111111111111111",
                "1111111111111111111111000111111111111111111110000111111111111111111111111111111111111111111111111111111110001111111111111111111100011111111111111111111111111111",
                "1111111111111111111111000111111111011111111110000111111111111111111111111111111111111111111111111111111110001111111111011111111100011111111111111111111111111111",
                "1111111111111111111111000111111110001111111110000111111111111111111111111111111111111111111111111111111110001111111110001111111100011111111111111111111111111111",
                "1111111111111111111111000111111100000111111110000111111111111111111111111111111111111111111111111111111110001111111100000111111100011111111111111111111111111111",
                "1111111111111111111111000111111000001111111110000111111111111111111111111111111111111111111111111111111110001111111110000011111100011111111111111111111111111111",
                "1111111111111111111111000111110000000001111110000111111111111111111111111111111111111111111111111111111110001111110000000001111100011111111111111111111111111111",
                "1111111111111111111111000111100000000000111110000111111111111111111111111111111111111111111111111111111110001111100000000000111100011111111111111111111111111111",
                "1111111111111111111111000111000000000000111110000111111111111111111111111111111111111111111111111111111110001111100000000000011100011111111111111111111111111111",
                "1111111111111111111111000111100000000000111110000111111111111111111111111111111111111111111111111111111110001111100000000000111100011111111111111111111111111111",
                "1111111111111111111111000111110000000001111110000111111111111111111111111111111111111111111111111111111110001111110000000001111100011111111111111111111111111111",
                "1111111111111111111111000111111000001111111110000111111111111111111111111111111111111111111111111111111110001111111110000011111100011111111111111111111111111111",
                "1111111111111111111111000111111100000111111110000111111111111111111111111111111111111111111111111111111110001111111100000111111100011111111111111111111111111111",
                "1111111111111111111111000111111110001111111110000111111111111111111111111111111111111111111111111111111110001111111110001111111100011111111111111111111111111111",
                "1111111111111111111111000111111111011111111110000111111111111111111111111111111111111111111111111111111110001111111111011111111100011111111111111111111111111111",
                "1111111111111111111111000111111111111111111110000111111111111111111111111111111111111111111111111111111110001111111111111111111100011111111111111111111111111111",
                "1111111111111111111111000111111111111111111110000111111111111111111111111111111111111111111111111111111110001111111111111111111100011111111111111111111111111111",
                "1111111111111111111111000111111111111111111110000111111111111111111111111111111111111111111111111111111110001111111111111111111100011111111111111111111111111111",
                "1111111111111111111111000000000000000000000000000111111111111111111111111111111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
                "1111111111111111111111000000000000000000000000001111111111111111111111111111111111111111111111111111111110000000000000000000000000011111111111111111111111111111",
                "1111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111",
                "1111111111111111111111110000000000000000000000111111111111111111111111111111111111111111111111111111111111100000000000000000000001111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111001111111111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111110000111111111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111110000111111111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111110010000100111111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111100000000000001111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111100000000000001111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111110000000000011111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111000000000111111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111100000001111111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111110000011111111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111000111111111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111101111111111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000111111111111111111111000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
                "1111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");
   
  BorderLine <=("000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",
                "011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110",                    
                "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000");

ArrowIngameLogoCircle <=
   ("11111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111",
    "11111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111",
    "11111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111",
    "11111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111",
    "11111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111",
    "11111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111",
    "11111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111",
    "11111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111",
    "11111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111",
    "11111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111",
    "11111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111",
    "11111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111",
    "11111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111",
    "11111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111",
    "11111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111",
    "11111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111",
    "11111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111",
    "11111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111",
    "11111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111",
    "11111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111",
    "11111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111",
    "11111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111",
    "11111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111",
    "11111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111",
    "11111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111",
    "11111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111",
    "11111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111",
    "11111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111",
    "11111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111",
    "11111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111",
    "11111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
    "11111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111",
    "11111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111",
    "11111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111",
    "11111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111",
    "11111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111",
    "11111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111",
    "11111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111",
    "11111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111",
    "11111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000111111000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111",
    "11111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111",
    "11111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111",
    "11111111111111000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111111",
    "11111111111111000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111111",
    "11111111111110000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111111",
    "11111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111111",
    "11111111111100000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111",
    "11111111111000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111111",
    "11111111110000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111",
    "11111111110000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000111111111",
    "11111111100000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000111111111",
    "11111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000011111111",
    "11111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000011111111",
    "11111111000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000001111111",
    "11111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000001111111",
    "11111110000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000111111",
    "11111100000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000111111",
    "11111100000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000111111",
    "11111100000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000011111",
    "11111000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000011111",
    "11111000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000001111",
    "11110000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000001111",
    "11110000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000001111",
    "11110000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000111",
    "11100000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000111",
    "11100000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000111",
    "11100000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000111",
    "11100000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000011",
    "11000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000011",
    "11000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000011",
    "11000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000011",
    "11000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000001",
    "11000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000001",
    "10000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000001",
    "10000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000001",
    "10000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000001",
    "10000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000",
    "00000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000",
    "10000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000",
    "10000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000",
    "10000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000",
    "11000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000",
    "11000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000",
    "11000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
    "11000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000",
    "11100000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000001",
    "11100000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000001",
    "11100000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000001",
    "11100000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000001",
    "11110000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000011",
    "11110000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000011",
    "11110000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000111",
    "11111000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000001111",
    "11111000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000001111",
    "11111000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000011111",
    "11111100000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000011111", 
    "11111100000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000011111", 
    "11111100000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000111111", 
    "11111110000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000111111", 
    "11111110000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000001111111", 
    "11111111000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000001111111", 
    "11111111000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000011111111", 
    "11111111100000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000011111111", 
    "11111111100000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000111111111", 
    "11111111110000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000111111111", 
    "11111111110000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111", 
    "11111111111000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000001111111111", 
    "11111111111000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000011111111111", 
    "11111111111100000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000111111111111", 
    "11111111111100000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000111111111111", 
    "11111111111110000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111111", 
    "11111111111111000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000011111111111111", 
    "11111111111111100000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111", 
    "11111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111", 
    "11111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000011111110000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111", 
    "11111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111", 
    "11111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111", 
    "11111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111", 
    "11111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111", 
    "11111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111", 
    "11111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111", 
    "11111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111", 
    "11111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111", 
    "11111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111", 
    "11111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111", 
    "11111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111", 
    "11111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111", 
    "11111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111", 
    "11111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111", 
    "11111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111", 
    "11111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111", 
    "11111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111", 
    "11111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111", 
    "11111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111", 
    "11111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111", 
    "11111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"); 
                                                                                                                                                                                                                                                                                                                                                                                                  
 ArrowInGameLogoArrow <=
   ("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111100000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111100000000000000000000000000000000010000000000000000000000010000000000000000000000000000000001111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111100000000000000000000000000000000110000000000000000000000011000000000000000000000000000000001111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111000000000000000000000000000000001110000000000000000000000011100000000000000000000000000000001111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111000000000000000000000000000000011110000000000000000000000011110000000000000000000000000000000111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111000000000000000000000000000000111110000000000000000000000011111000000000000000000000000000000111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111000000000000000000000000000001111110000000000000000000000011111100000000000000000000000000000111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111000000000000000000000000000011111110000000000000000000000011111110000000000000000000000000000111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111000000000000000000000000000111111110000000000000000000000011111111000000000000000000000000000111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111000000000000000000000000001111111110000000000000000000000011111111100000000000000000000000001111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111100000000000000000000000011111111110000000000000000000000011111111110000000000000000000000001111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111100000000000000000000000111111111110000000000000000000000011111111111000000000000000000000001111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111110000000000000000000001111111111110000000000000000000000011111111111100000000000000000000011111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111000000000000000000011111111111110000000000000000000000011111111111110000000000000000000111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111100000000000000000111111111111110000000000000000000000011111111111111000000000000000001111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111110000000000000001111111111111110000000000000000000000011111111111111100000000000000011111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111000000000000011111111111111110000000000000000000000011111111111111110000000000000111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111100000000000111111111111111110000000000000000000000011111111111111111000000000001111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111110000000001111111111111111110000000000000000000000011111111111111111100000000011111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111100000111111111111111111110000000000000000000000011111111111111111111000001111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",                                                                                                                                                                                                             
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",  
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",  
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",  
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",  
    "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111"); 
    
    
 ARRHYTHMIA_IN_GAME <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111110000000000000000011111111100000000000000000001111111111110000000000000000001111111111110000000011110000000000111110000000000000000000000011110000000000000000000000011111000000000000110000000000001111110000000000011100000000000111100000000000011111111110000000000000000000011111111111111",
"111111111111100000000000000000000111110000000000000000000000001111111000000000000000000000001111111000000000000110000000000001110000000000000000000000011110000000000000000000000001111000000000000110000000000001111100000000000001000000000000111100000000000001111111110000000000000000000011111111111111",
"111111111111000000000000000000000111110000000000000000000000001111111000000000000000000000001111111000000000000100000000000001110000000000000000000000011110000000000000000000000001111000000000000010000000000001111100000000000011000000000000111100000000000001111111110000000000000000000011111111111111",
"111111111111100000000000000000000111110000000000000000000000001111111000000000000000000000001111111000000000000100000000000001110000000000000000000000011110000000000000000000000001111000000000000010000000000001111100000000000011000000000000111100000000000001111111110000000000000000000011111111111111",
"111111111111000000000000000000000111110000000000000000000000001111111000000000000000000000001111111000000000000100000000000001110000000000000000000000000110000000000000000000000000111000000000000000000000000000011100000000000000000000000000011100000000000000111110000000000000000000000001111111111111",
"111111111100000000000000000000000001110000000000000000000000000011111000000000000000000000000011111000000000000000000000000000110000000000000000000000000010000000000000000000000000011000000100000000000000000000001100000000000000000000000000001100000000000000011100000000000000000000000000011111111111",
"111111111000000011111111111100000000110000011111111111111000000011111000011111111111111100000011111000001110000000000111100000010000111100000001111000000010000011111111111111000000011000001110000000000111110000001100000111100000000011110000000100000111100000011100000001111111111110000000011111111111",
"111111111000000011111111111100000000110000011111111111111100000011111000011111111111111100000011111000001110000000000111100000010000111100000001111000000010000011111111111111000000011000001110000000000111100000001100000111100000000001110000000100000111100000011100000001111111111110000000011111111111",
"111111111000000011111111111100000000110000011111111111111100000011111000011111111111111100000011111000001110000000000111100000010000111100000001111000000010000000011111110000000000011000001110000000000111100000001100000111100000000011110000000100000111000000011100000001110000000110000000001111111111",
"111111111000000011100000001110000000010000011110000000001100000000111000011111000000001100000000111000001110000000000111100000010000111100000001111000000010000000000111100000000000011000001110000000000111100000001100000111110000000111110000000100000111000000011100000011100000000011100000000111111111",
"111111111000001111000000000111100000010000011110000000000110000000111000011110000000000111000000011000001110000000000111100000010000111100000001111000000010000000000111000000000000011000001110000000000111100000001100000111111000001111110000000100000111000000011100000111100000000001110000000111111111",
"111111111000001111000000000011100000010000011100000000000111000000011000011110000000000111100000011000001110000000000111100000010000111100000001111000000010000000000111000000000000011000001110000000000111100000001100000111111000011111110000000100000111000000011100000111100000000001111000000111111111",
"111111111000001111000000000011100000010000011100000000000111000000011000011110000000000111100000011000001110000000000111100000010000111100000001111000000010000000000111000000000000011000001110000000000111100000001100000111111000011111110000000100000111000000011100000111100000000001111000000111111111",
"111111111000001111000000000011100000010000011100000000000111000000011000011110000000000111100000011000001110000000000111100000010000111100000001111000000011100000000111000000000000011000001110000000000111100000001100000111111111111111110000000100000111000000011100000111100000000001111000000111111111",
"111111111000001111000000000011100000010000011100000000000111000000011000011110000000000111100000011000001110000000000111100000010000111100000001111000000011111100000111000000000000011000001110000000000111100000001100000111111111111111110000000100000111000000011100000111100000000001111000000111111111",
"111111111000001111000000000011100000010000011100000000000111000000011000011110000000000111100000011000001110000000000111100000010000111100000001111000000011111100000111000000000000011000001110000000000111100000001100000111111111111111110000000100000111000000011100000111100000000001111000000111111111",
"111111111000001111000000000011100000010000011100000000000111000000011000011110000000000111100000011000001110000000000111100000010000111100000001110000000011111100000111000000000000011000001110000000000111100000001100000111111111111111110000000100000111000000011100000111100000000001111000000111111111",
"111111111000001111000000000011100000010000011110000000001100000000011000011110000000001110000000011000001110000000000111100000010000000110000011000000000011111100000111000000000000111000001111000000000111100000001100000111100001000011110000000100000111000000011100000111100000000001111000000111111111",
"111111111000001111000000000011100000010000011111100000111100000000011000011111100000111100000000011000001111111111111111100000010000000111111111000000000011111100000111000000011111111000001111111111111111100000001100000111000001000001110000000100000111000000011100000111100000000001111000000111111111",
"111111111000001111000000000011100000010000011111111111111100000000011000011111111111111100000000011000001111111111111111100000010000000111111111000000000011111100000111000000011111111000001111111111111111100000001100000111000001000001110000000100000111000000011100000111100000000001111000000111111111",
"111111111000001111000000000011100000010000011111111111111100000000011000011111111111111100000000011000001111111111111111100000010000000011111111000000000011111100000111000000001111111000001111100000001111100000001100000111100000000001110000000100000111000000011100000111100000000011111000000111111111",
"111111111000001111000000000111100000010000011100000000000100000000011000011111000000001100000000011000001111000000001111100000011000000001111100000000000011111100000111000000001111111000001110000000000111100000001100000111100000000001110000000100000111000000011100000111110000000111111000000111111111",
"111111111000001111111111111111100000010000011100000000000110000000011000011110000000000111000000011000001110000000000111100000001100000000111000000000000011111100000111000000001111111000001110000000000111100000001100000111100000000001110000000100000111000000011100000111111111111111111000000111111111",
"111111111000001111111111111111100000010000011100000000000111000000011000011110000000000111100000011000001110000000000111100000001110000000111000000000000011111100000111000000001111111000001110000000000111100000001100000111100000000001110000000100000111000000011100000111111111111111111000000111111111",
"111111111000001111111111111111100000010000011100000000000111000000011000011110000000000111100000011000001110000000000111100000001110000000111000000000000011111100000111000000001111111000001110000000000111100000001100000111100000000001110000000100000111000000011100000111111111111111111000000111111111",
"111111111000001111111111111111100000010000011100000000000111000000011000011110000000000111100000011000001110000000000111100000001110000000111000000000000011111100000111000000001111111000001110000000000111100000001100000111100000000001110000000100000111000000011100000111100000000011111000000111111111",
"111111111000001111000000000111100000010000011100000000000111000000011000011110000000000111100000011000001110000000000111100000001111000000111000000000001111111100000111000000001111111000001110000000000111100000001100000111100000000001110000000100000111000000011100000111100000000001111000000111111111",
"111111111000001111000000000011100000010000011100000000000111000000011000011110000000000111100000011000001110000000000111100000001111100000111000000000011111111100000111000000001111111000001110000000000111100000001100000111100000000001110000000100000111000000011100000111100000000001111000000111111111",
"111111111000001111000000000011100000010000011100000000000111000000011000011110000000000111100000011000001110000000000111100000001111100000111000000000011111111100000111000000001111111000001110000000000111100000001100000111100000000001110000000100000111000000011100000111100000000001111000000111111111",
"111111111000001111000000000011100000010000011100000000000111000000011000011110000000000111100000011000001110000000000111100000001111100000111000000000111111111100000111000000001111111000001110000000000111100000001100000111100000000001110000000100000111000000011100000111100000000001111000000111111111",
"111111111000001111000000000011100000010000011100000000000111000000011000011110000000000111100000011000001110000000000111100000001111100000111000000001111111111100000111000000001111111000001110000000000111100000001100000111100000000001110000000100000111000000011100000111100000000001111000000111111111",
"111111111000001111000000000011100000010000011100000000000111000000011000011110000000000111100000011000001110000000000111100000001111100000111000000011111111111100000111000000001111111000001110000000000111100000001100000111100000000011110000000100000111100000011100000111100000000011111000000111111111",
"111111111000001111000000000111100000010000011100000000000111000000011000011110000000000111100000011000001110000000000111100000001111100000111000000001111111111100000111000000001111111000001110000000000111100000001100000111100000000011110000000100000111100000011100000111100000000011111000000111111111",
"111111111000001111000000000011100000010000011100000000000111000000011000001110000000000111100000011000001110000000000111100000001111100000000000000001111111111100000010000000001111111000000100000000000000000000001100000001000000000000100000000100000000000000011100000000000000000000000000000111111111",
"111111111000000000000000000000000000010000000000000000000000000000011000000000000000000000000000011000000000000000000000000000001111100000000000000001111111111100000000000000001111111000000000000000000000000000001100000000000000000000000000000100000000000000011100000000000000000000000000000111111111",
"111111111000000000000000000000000000010000000000000000000000000000011000000000000000000000000000011000000000000000000000000000001111100000000000000001111111111100000000000000001111111000000000000000000000000000001100000000000000000000000000000100000000000000011100000000000000000000000000000111111111",
"111111111000000000000000000000000000010000000000000000000000000000011000000000000000000000000000011000000000000000000000000000001111100000000000000001111111111100000000000000001111111000000000000000000000000000001100000000000000000000000000000100000000000000011100000000000000000000000000000111111111",
"111111111000000000000000000000000000010000000000000000000000000000011000000000000000000000000000011000000000000000000000000000001111100000000000000001111111111110000000000000001111111000000000000000000000000000001110000000000000000000000000000100000000000000011100000000000000000000000000000111111111",
"111111111000000000000000000000000000010000000000000000000000000000011000000000000000000000000000011000000000000000000000000000001111111000000000000001111111111111000000000000001111111100000000000000000000000000001111000000000000000000000000000111000000000000011110000000000000000000000000000111111111",
"111111111111000000000000000000000000011110000000000001100000000000011110000000000000100000000000011110000000000000100000000000001111111100000000000001111111111111100000000000001111111111000000000000110000000000001111100000000000011000000000000111100000000000011111110000000000011000000000000111111111",
"111111111111000000000000110000000000011110000000000001100000000000011110000000000001110000000000001111000000000001110000000000001111111100000000000001111111111111100000000000001111111111000000000000110000000000001111100000000000011000000000000111100000000000011111110000000000011000000000000111111111",
"111111111111000000000000110000000000011110000000000001100000000000011110000000000001110000000000001111000000000001110000000000001111111100000000000011111111111111100000000000001111111111000000000000110000000000001111100000000000011000000000000111100000000000011111110000000000011000000000000111111111",
"111111111111100000000000110000000000011110000000000001100000000000011110000000000001110000000000011111000000000001110000000000011111111110000000000011111111111111110000000000011111111111100000000001111000000000011111110000000000011100000000001111110000000000011111110000000000011100000000000111111111",
"111111111111110000000111111110000000111111110000000111111000000001111111110000000111111000000001111111110000000111111100000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
"111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");
   
    
    
    
    
 UP_Arrow <= 
              ("11111111111111111111111111111111111111111111111111",
               "11111111111111111111111100111111111111111111111111",
               "11111111111111111111111000011111111111111111111111",
               "11111111111111111111111000011111111111111111111111",
               "11111111111111111111110000001111111111111111111111",
               "11111111111111111111100000000111111111111111111111",
               "11111111111111111111100000000111111111111111111111",
               "11111111111111111111000000000011111111111111111111",
               "11111111111111111110000011000001111111111111111111",
               "11111111111111111110000011000001111111111111111111",
               "11111111111111111100000111100000111111111111111111",
               "11111111111111111000001111110000011111111111111111",
               "11111111111111110000001111110000001111111111111111",
               "11111111111111110000011111111000001111111111111111",
               "11111111111111100000111111111100000111111111111111",
               "11111111111111000000111111111100000011111111111111",
               "11111111111111000001111111111110000011111111111111",
               "11111111111110000011111100111111000001111111111111",
               "11111111111100000011111000011111000000111111111111",
               "11111111111100000111110011001111100000111111111111",
               "11111111111000001111000111100011110000011111111111",
               "11111111110000001111000111100011110000001111111111",
               "11111111110000011110000111100001111000001111111111",
               "11111111100000111100000111100000111100000111111111",
               "11111111000001111100000111100000111110000011111111",
               "11111111000001111000000111100000011110000011111111",
               "11111111000001110000000111100000001110000011111111",
               "11111111000001100000000111100000000110000011111111",
               "11111111000000000000000100100000000000000011111111",
               "11111111000000000000000000000000000000000011111111",
               "11111111000000000000000011000000000000000011111111",
               "11111111100000000000000111100000000000000111111111",
               "11111111100000000110000111100001100000000111111111",
               "11111111110000001110000111100001110000001111111111",
               "11111111111000001110000111100001110000011111111111",
               "11111111111110111110000111100001111101111111111111",
               "11111111111111111110000111100001111111111111111111",
               "11111111111111111110000111100001111111111111111111",
               "11111111111111111110000111100001111111111111111111",
               "11111111111111111110000111100001111111111111111111",
               "11111111111111111110000011000001111111111111111111",
               "11111111111111111110000000000001111111111111111111",
               "11111111111111111110000000000001111111111111111111",
               "11111111111111111111000000000011111111111111111111",
               "11111111111111111111100000000111111111111111111111",
               "11111111111111111111100000000111111111111111111111",
               "11111111111111111111110000001111111111111111111111",
               "11111111111111111111111000011111111111111111111111",
               "11111111111111111111111000111111111111111111111111",
               "11111111111111111111111100111111111111111111111111");

 Down_Arrow <= 
               ("11111111111111111111111100111111111111111111111111",
                "11111111111111111111111100011111111111111111111111",
                "11111111111111111111111000011111111111111111111111",
                "11111111111111111111110000001111111111111111111111",
                "11111111111111111111100000000111111111111111111111",
                "11111111111111111111100000000111111111111111111111",
                "11111111111111111111000000000011111111111111111111",
                "11111111111111111110000000000001111111111111111111",
                "11111111111111111110000000000001111111111111111111",
                "11111111111111111110000011000001111111111111111111",
                "11111111111111111110000111100001111111111111111111",
                "11111111111111111110000111100001111111111111111111",
                "11111111111111111110000111100001111111111111111111",
                "11111111111111111110000111100001111111111111111111",
                "11111111111110111110000111100001111101111111111111",
                "11111111111000001110000111100001110000011111111111",
                "11111111110000001110000111100001110000001111111111",
                "11111111100000000110000111100001100000000111111111",
                "11111111100000000000000111100000000000000111111111",
                "11111111000000000000000011000000000000000011111111",
                "11111111000000000000000000000000000000000011111111",
                "11111111000000000000000100100000000000000011111111",
                "11111111000001100000000111100000000110000011111111",
                "11111111000001110000000111100000001110000011111111",
                "11111111000001111000000111100000011110000011111111",
                "11111111000001111100000111100000111110000011111111",
                "11111111100000111100000111100000111100000111111111",
                "11111111110000011110000111100001111000001111111111",
                "11111111110000001111000111100011110000001111111111",
                "11111111111000001111000111100011110000011111111111",
                "11111111111100000111110011001111100000111111111111",
                "11111111111100000011111000011111000000111111111111",
                "11111111111110000011111100111111000001111111111111",
                "11111111111111000001111111111110000011111111111111",
                "11111111111111000000111111111100000011111111111111",
                "11111111111111100000111111111100000111111111111111",
                "11111111111111110000011111111000001111111111111111",
                "11111111111111110000001111110000001111111111111111",
                "11111111111111111000001111110000011111111111111111",
                "11111111111111111100000111100000111111111111111111",
                "11111111111111111110000011000001111111111111111111",
                "11111111111111111110000011000001111111111111111111",
                "11111111111111111111000000000011111111111111111111",
                "11111111111111111111100000000111111111111111111111",
                "11111111111111111111100000000111111111111111111111",
                "11111111111111111111110000001111111111111111111111",
                "11111111111111111111111000011111111111111111111111",
                "11111111111111111111111000011111111111111111111111",
                "11111111111111111111111100111111111111111111111111",
                "11111111111111111111111111111111111111111111111111");
            
 Left_Arrow <=
               ("11111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111",
                "11111111111111111111111100000001111111111111111111",
                "11111111111111111111111000000000011111111111111111",
                "11111111111111111111100000000000001111111111111111",
                "11111111111111111111000000000000000111111111111111",
                "11111111111111111100000000000000000111111111111111",
                "11111111111111111000000011110000000011111111111111",
                "11111111111111100000000111110000000111111111111111",
                "11111111111111000000001111100000000111111111111111",
                "11111111111100000000111111000000011111111111111111",
                "11111111111000000001111110000000111111111111111111",
                "11111111110000000111111000000000111111111111111111",
                "11111111000000001111110000000000000000000001111111",
                "11111110000000111111000000000000000000000000111111",
                "11111000000001111111000000000000000000000000001111",
                "11110000000111111110000000000000000000000000000111",
                "11000000001111111100111111111001111111110000000011",
                "10000000111111111001111111110011111111111000000000",
                "10000000111111111001111111110011111111111000000000",
                "11000000001111111100111111111001111111110000000001",
                "11110000000111111110000000000000000000000000000111",
                "11111000000001111111000000000000000000000000001111",
                "11111110000000111111000000000000000000000000111111",
                "11111111000000001111110000000000000000000001111111",
                "11111111110000000111111000000000111111111111111111",
                "11111111111000000001111110000000111111111111111111",
                "11111111111100000000111111000000011111111111111111",
                "11111111111111000000001111100000000111111111111111",
                "11111111111111100000000111110000000111111111111111",
                "11111111111111111000000011110000000011111111111111",
                "11111111111111111100000000000000000111111111111111",
                "11111111111111111111000000000000000111111111111111",
                "11111111111111111111100000000000001111111111111111",
                "11111111111111111111111000000000011111111111111111",
                "11111111111111111111111100000001111111111111111111",
                "11111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111",
                "11111111111111111111111111111111111111111111111111");
        
 Right_Arrow  <=
              ("11111111111111111111111111111111111111111111111111",  
               "11111111111111111111111111111111111111111111111111",  
               "11111111111111111111111111111111111111111111111111",  
               "11111111111111111111111111111111111111111111111111",  
               "11111111111111111111111111111111111111111111111111",  
               "11111111111111111111111111111111111111111111111111",  
               "11111111111111111111111111111111111111111111111111",  
               "11111111111111111111111111111111111111111111111111",  
               "11111111111111111110000000111111111111111111111111",  
               "11111111111111111000000000011111111111111111111111",  
               "11111111111111110000000000000111111111111111111111",  
               "11111111111111100000000000000011111111111111111111",  
               "11111111111111100000000000000000111111111111111111",  
               "11111111111111000000001111000000011111111111111111",  
               "11111111111111100000001111100000000111111111111111",  
               "11111111111111100000000111110000000011111111111111",  
               "11111111111111111000000011111100000000111111111111",  
               "11111111111111111100000001111110000000011111111111",  
               "11111111111111111100000000011111100000001111111111",  
               "11111110000000000000000000001111110000000011111111",  
               "11111100000000000000000000000011111100000001111111",  
               "11110000000000000000000000000011111110000000011111",  
               "11100000000000000000000000000001111111100000001111",  
               "10000000001111111110011111111100111111110000000011",  
               "00000000011111111111001111111110011111111100000001",  
               "00000000011111111111001111111110011111111100000001",  
               "11000000001111111110011111111100111111110000000011",  
               "11100000000000000000000000000001111111100000001111",  
               "11110000000000000000000000000011111110000000011111",  
               "11111100000000000000000000000011111100000001111111",  
               "11111110000000000000000000001111110000000011111111",  
               "11111111111111111100000000011111100000001111111111",  
               "11111111111111111100000001111110000000011111111111",  
               "11111111111111111000000011111100000000111111111111",  
               "11111111111111100000000111110000000011111111111111",  
               "11111111111111100000001111100000000111111111111111",  
               "11111111111111000000001111000000011111111111111111",  
               "11111111111111100000000000000000111111111111111111",  
               "11111111111111100000000000000011111111111111111111",  
               "11111111111111110000000000000111111111111111111111",  
               "11111111111111111000000000011111111111111111111111",  
               "11111111111111111110000000111111111111111111111111",  
               "11111111111111111111111111111111111111111111111111",  
               "11111111111111111111111111111111111111111111111111",  
               "11111111111111111111111111111111111111111111111111",  
               "11111111111111111111111111111111111111111111111111",  
               "11111111111111111111111111111111111111111111111111",  
               "11111111111111111111111111111111111111111111111111",  
               "11111111111111111111111111111111111111111111111111",  
               "11111111111111111111111111111111111111111111111111"); 
               

PERFECT<=
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000011111111000000000000000001111111000000000000000000000111111",
 "11111111111111111111111111111111000000000000000000000000111110000000000000000000001111111100000000000000000000000111100000000000000000000000011111110000000000000000001111111000000000000000000000111111",
 "11110000000000000000000001111111000000000000000000000000111110000000000000000000001111111100000000000000000000000111100000000000000000000000011111110000000000000000001111111000000000000000000000111111",
 "11110000000000000000000011111111000000000000000000000000111110000000000000000000001111111100000000000000000000000111100000000000000000000000011111110000000000000000001111111000000000000000000000111111",
 "11110000000000000000000011111111000000000000000000000000111110000000000000000000001111111100000000000000000000000111100000000000000000000000011111110000000000000000001111111000111111111111111000111111",
 "11110000000000000000000011111111000000000000000000000000111110000000000000000000001111111100000000000000000000000111100011111111111111111100000111000001111111111111000001111000111111111111111100000111",
 "11110001111111111111110001111111000111111111111111111000001110001111111111111111000001111100111111111111111111100001100011111111111111111100000111000001111111111111000001111000111111111111111100000111",
 "11110011111111111111110000011111000111111111111111111000001110001111111111111111000001111100111111111111111111100001100011111111111111111100000111000001111111111111000001111000111111111111111100000111",
 "11110011111111111111110000011111000111111111111111111000001110001111111111111111000001111100111111111111111111100001100011111111111111111100000111000001111111111111000001111000111111111111111100000111",
 "11110011111111111111110000011111000111111111111111111000001110001111111111111110000001111100111111111111111111100001100011111111111111111100000111000001111111111111000001111000000001111100000000000111",
 "11110011111111111111110000011111000111111111111111111000001110001111111111111111110001111100111111111111111111000001100011111000000000000000000111001111110000000111111000011000000001111100000000000111",
 "11110011111100000001111110010111000111110000000000000000001110001111100000000111110000011100111111000000000000000001100011111000000000000000000111001111110000000111111000011000000001111100000000000111",
 "11110011111100000001111110000111000111110000000000000000001110001111100000000111110000011100111111000000000000000001100011111000000000000000000111001111110000000111111000011000000001111100000000000111",
 "11110011111100000001111110000111000111110000000000000000001110001111100000000111110000011100111111000000000000000001100011111000000000000000000111001111110000000111111000011111111001111100000000000111",
 "11110011111100000001111110000111000111110000000000000000001110001111100000000111110000011100111111000000000000000001100011111000000000000000000111001111110000000000000000011111111001111100000000000111",
 "11110011111100000001111110000111000111110000000000000000001110001111100000000111110000011100111111000000000000000001100011111000000000000000000111001111110000000000000000011111111001111100000000000111",
 "11110011111100000001111110000111000111110000000000000000001110001111100000000111110000011100111111000000000000000001100011111000000000000000000111001111110000000000000000011111111001111100000000000111",
 "11110011111100000001111110000111000111110000000000000000001110001111100000000111110000011100111111000000000000000001100011111000000000000000000111001111110000000000000000011111111001111100000000000111",
 "11110011111100000001111110000111000111110000000000000000001110001111100000000111110000011100111111000000000000000001100011111100000000000000000111001111110000000000000000011111111001111100000111111111",
 "11110011111100000001111110000111000111111111111111000000111110001111111111111111110000011100111111111111111100000111100011111111111111110000011111001111110000000000000000011111111001111100000111111111",
 "11110011111100000001111110000111000111111111111111100000111110001111111111111110000000011100111111111111111100000111100011111111111111110000011111001111110000000000000000011111111001111100000111111111",
 "11110011111100000001111110000111000111111111111111000000111110001111111111111111000000011100111111111111111100000111100011111111111111110000011111001111110000000000000000011111111001111100000111111111",
 "11110011111100000001111110000111000111111111111111000000111110001111111111111110000000011100111111111111111100000111100011111111111111110000011111001111110000000000000000011111111001111100000111111111",
 "11110011111100000001111110000111000111111111111111000000111110001111111111111111000000011100111111111111111100000111100011111100000000000000011111001111110000000000000001111111111001111100000111111111",
 "11110011111111111111111100000111000111110000000000000000111110001111100000000111110000011100111111000000000000000111100011111000000000000000011111001111110000000000000001111111111001111100000111111111",
 "11110011111111111111110000000111000111110000000000000000111110001111100000000111110000011100111111000000000000000111100011111000000000000000011111001111110000000000000001111111111001111100000111111111",
 "11110011111111111111110000000111000111110000000000000000111110001111100000000111110000011100111111000000000000000111100011111000000000000000011111001111110000000000000001111111111001111100000111111111",
 "11110011111111111111110000000111000111110000000000000000111110001111100000000111110000011100111111000000000000000111100011111000000000000000011111001111110000000000000001111111111001111100000111111111",
 "11110011111111111111110000000111000111110000000000000000111110001111100000000111110000011100111111000000000000000111100011111000000000000000011111001111110000000111111000011111111001111100000111111111",
 "11110011111111111111110000000111000111110000000000000000111110001111100000000111110000011100111111000000000000000111100011111000000000000000011111001111110000000111111000011111111001111100000111111111",
 "11110011111100000000000000000111000111110000000000000000111110001111100000000111110000011100111111000000000000000111100011111000000000000000011111001111110000000111111000011111111001111100000111111111",
 "11110011111100000000000000000111000111110000000000000000111110001111100000000111110000011100111111000000000000000111100011111000000000000000011111001111110000000111111000011111111001111100000111111111",
 "11110011111100000000000000000111000111110000000000000000111110001111100000000111110000011100111111000000000000000111100011111111111111111100000111001111111111111111111000011111111001111100000111111111",
 "11110011111100000000000000000111000111111111111111111000001110001111100000000111110000011100111111000011111111111111100011111111111111111100000111000001111111111111000000011111111001111100000111111111",
 "11110011111100000000000000011111000111111111111111111000001110001111100000000111110000011100111111000011111111111111100011111111111111111100000111000001111111111111000000011111111001111100000111111111",
 "11110011111100000000000000011111000111111111111111111000001110001111100000000111110000011100111111000011111111111111100011111111111111111100000111000001111111111111000000011111111001111100000111111111",
 "11110011111100000000000000011111000111111111111111111000001110001111100000000111110000011100111111000011111111111111100011111111111111111100000111000001111111111111000000011111111001111100000111111111",
 "11110011111100000000000000011111000111111111111111111000001110001111100000000111110000011100111111000011111111111111100011111111111111111100000111110001111111111111000000011111111000000000000111111111",
 "11110011111100000000000000011111000111111111111111111000001110000000000000000000000000011100000000000011111111111111100000000000000000000000000111110000000000000000000000011111111000000000000111111111",
 "11110000000000001111111111111111000000000000000000000000001110000000000000000000000000011100000000000011111111111111100000000000000000000000000111110000000000000000000000011111111000000000000111111111",
 "11110000000000001111111111111111000000000000000000000000001110000000000000000000000000011100000000000011111111111111100000000000000000000000000111110000000000000000000000011111111000000000000111111111",
 "11110000000000001111111111111111000000000000000000000000001110000000000000000000000000011100000000000011111111111111110000000000000000000000000111111000000000000000000000011111111110000000000111111111",
 "11110000000000001111111111111111111000000000000000000000001111110000000000111000000000011111000000000011111111111111111100000000000000000000000111111110000000000000000001111111111111000000000111111111",
 "11111100000000001111111111111111111000000000000000000000001111110000000000111000000000011111000000000011111111111111111100000000000000000000000111111110000000000000000001111111111111000000000111111111",
 "11111110000000001111111111111111111000000000000000000000001111110000000000111000000000011111000000000011111111111111111100000000000000000000000111111110000000000000000001111111111110000000000111111111",
 "11111110000000001111111111111111111000000000000000000000001111110000000000111000000000011111000000000011111111111111111100000000000000000000000111111110000000000000000001111111111111000000000111111111",
 "11111110000000001111111111111111111000000000000000000000001111110000000000111000000000011111000000000011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111110000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



GOOD   <=
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111110000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111110000000000000000000000000000001111111111111111110000000000000000000000000000001111111111111111110000000000000000000000000000001111111111110000000000000000000000000000001111111111111111111",
 "11111111111110000000000000000000000000000001111111111111111110000000000000000000000000000001111111111111111110000000000000000000000000000001111111111110000000000000000000000000000001111111111111111111",
 "11111111111110000000000000000000000000000001111111111111111110000000000000000000000000000001111111111111111110000000000000000000000000000001111111111110000000000000000000000000000001111111111111111111",
 "11111111111110000000000000000000000000000001111111111111111110000000000000000000000000000001111111111111111110000000000000000000000000000001111111111110000000000000000000000000000001111111111111111111",
 "11111111000000000111111111111111111111100000000111111111111100000111111111111111111111000001111111111111111100000111111111111111111111000001111111111110000011111111111111111111100001111111111111111111",
 "11111111000000000111111111111111111111100000000111111111000000001111111111111111111111000000000111111111000000001111111111111111111111000000000111111110000111111111111111111111100000000011111111111111",
 "11111111000000000111111111111111111111100000000111111111000000001111111111111111111111000000000111111111000000001111111111111111111111000000000111111110000111111111111111111111100000000011111111111111",
 "11111111000000000111111111111111111111100000000111111111000000001111111111111111111111000000000111111111000000001111111111111111111111000000000111111110000111111111111111111111100000000011111111111111",
 "11111111000001111111110000000000001111111110000000011111000000001111111111111111111111100000000111111111000000001111111111111111111111100000000111111110000111111111111111111111110000000011111111111111",
 "11111111000001111111110000000000001111111110000000011111000011111111110000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000001111111110000000001111111111",
 "11111111000001111111110000000000001111111110000000011111000011111111100000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000001111111110000000001111111111",
 "11111111000001111111110000000000001111111110000000011111000011111111100000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000001111111110000000001111111111",
 "11111111000001111111110000000000000000000000000000011111000011111111100000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000001111111111001000001111111111",
 "11111111000001111111110000000000000000000000000000011111000011111111100000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000000000011111111100000000111111",
 "11111111000001111111110000000000000000000000000000011111000011111111100000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000000000011111111100000000111111",
 "11111111000001111111110000000000000000000000000000011111000011111111100000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000000000011111111100000000111111",
 "11111111000001111111110000000011111111111110000000011111000011111111100000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000000000011111111100000000111111",
 "11111111000001111111110000000111111111111110000000011111000011111111100000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000000000011111111100000000111111",
 "11111111000001111111110000000111111111111110000000011111000011111111100000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000000000011111111100000000111111",
 "11111111000001111111110000000111111111111110000000011111000011111111100000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000000000011111111100000000111111",
 "11111111000001111111110000000011101111111110000000011111000011111111100000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000000000011111111100000000111111",
 "11111111000001111111110000000000001111111110000000011111000011111111100000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000000000011111111100000000111111",
 "11111111000001111111110000000000001111111110000000011111000011111111100000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000000000011111111100000000111111",
 "11111111000001111111110000000000001111111110000000011111000011111111100000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000000000011111111100000000111111",
 "11111111000001111111110000000000001111111110000000011111000011111111100000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000000000011111111100000000111111",
 "11111111000001111111110000000000001111111110000000011111000011111111100000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000000110111111111100000000111111",
 "11111111000001111111110000000000001111111110000000011111000011111111100000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000001111111110000000000000111111",
 "11111111000001111111110000000000001111111110000000011111000011111111100000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000001111111110000000000000111111",
 "11111111000001111111110000000000001111111110000000011111000011111111100000000000001111111110000000011111000011111111100000000000001111111110000000011110000111111111000000001111111110000000000000111111",
 "11111111000000000111111111111111110000111110000000011111000001111111110111111111111111111110000000011111000011111111111111111111111111111110000000011110000111111111100000001111111110000000000000111111",
 "11111111000000000111111111111111110000111110000000011111000000001111111111111111111111000000000000011111000000001111111111111111111111000000000000011110000111111111111111111111100000000000000000111111",
 "11111111000000000111111111111111110000111110000000011111000000001111111111111111111111000000000000011111000000001111111111111111111111000000000000011110000111111111111111111111100000000000000000111111",
 "11111111000000000111111111111111111000111110000000011111000000001111111111111111111111000000000000011111000000001111111111111111111111000000000000011110000111111111111111111111100000000000000000111111",
 "11111111100000000111111111111111110000111110000000011111000000001111111111111111111111000000000000011111000000001111111111111111111111000000000000011110000111111111111111111111100000000000000000111111",
 "11111111111110000000000000000000000000000000000000011111111100000111111111111111111111000000000000011111111100000111111111111111111111000000000000011110000011111111111111111111100000000000001111111111",
 "11111111111110000000000000000000000000000000000000011111111110000000000000000000000000000000000000011111111110000000000000000000000000000000000000011110000000000000000000000000000000000000001111111111",
 "11111111111110000000000000000000000000000000000000011111111110000000000000000000000000000000000000011111111110000000000000000000000000000000000000011110000000000000000000000000000000000000001111111111",
 "11111111111110000000000000000000000000000000000000011111111110000000000000000000000000000000000000011111111110000000000000000000000000000000000000011110000000000000000000000000000000000000001111111111",
 "11111111111111111000000000000000000000000000000000011111111111111000000000000000000000000000000111111111111111110000000000000000000000000000000111111111111000000000000000000000000000000011111111111111",
 "11111111111111111000000000000000000000000000000000011111111111111000000000000000000000000000000111111111111111111000000000000000000000000000000111111111111100000000000000000000000000000011111111111111",
 "11111111111111111000000000000000000000000000000000011111111111111000000000000000000000000000000111111111111111111000000000000000000000000000000111111111111100000000000000000000000000000011111111111111",
 "11111111111111111000000000000000000000000000000000011111111111111000000000000000000000000000000111111111111111111000000000000000000000000000000111111111111100000000000000000000000000000011111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111000000000000000000000000000001111111111111111111000000000000000000000000000001111111111111100000000000000000000000000000111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");







GREAT  <=
("11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111100000000000000000000000001111111111100000000000000000000000000001111111111100000000000000000000000000000000111111111110000000000000000000000000111111111100000000000000000000000000000111111111",
 "11111111100000000000000000000000001111111111100000000000000000000000000001111111111100000000000000000000000000000000111111111110000000000000000000000000111111111100000000000000000000000000000111111111",
 "11111111100000000000000000000000001111111111100000000000000000000000000001111111111100000000000000000000000000000000111111111110000000000000000000000000111111111100000000000000000000000000000111111111",
 "11111111100000000000000000000000001111111111100000000000000000000000000001111111111100000000000000000000000000000000111111111110000000000000000000000000111111111100000000000000000000000000000111111111",
 "11111111100000000000000000000000001111111111100000000000000000000000000001111111111100000000000000000000000000000000111111110000001111111111111111110000000111111100001111111111111111111110000000111111",
 "11111000000011111111111111111100000001111111100011111111111111111111110000001111111100001111111111111111111111111000000111100000001111111111111111110000000111111100001111111111111111111110000000011111",
 "11111000000011111111111111111100000001111111100011111111111111111111110000000111111100001111111111111111111111111000000111100000001111111111111111110000000111111100001111111111111111111110000000111111",
 "11111000000011111111111111111100000001111111100011111111111111111111110000000111111100001111111111111111111111111000000111100000001111111111111111110000000111111100001111111111111111111110000000111111",
 "11111000000011111111111111111100000001111111100011111111111111111111110000001111111100001111111111111111111111111000000111100000111111111111111111111111000011111100001111111111111111111110000000111111",
 "11111000011111111111111111111111110001111111100011111111111111111111111110000111111100001111111111111111111111111000000111100001111111100000000001111111000000011100000000000111111100000000000000111111",
 "11111000011111110000000000011111110000001111100011111111000000000011111110000000111100001111111000000000000000000000000111100001111111100000000001111111000000011100000000000111111100000000000000111111",
 "11111000011111110000000000011111110000001111100011111111000000000011111110000000111100001111111000000000000000000000000111100001111111100000000001111111000000011100000000000111111100000000000000111111",
 "11111000011111110000000000111111110000001111100011111111000000000011111110000000111100001111111000000000000000000000000111100001111111100000000001111111000000011110000000000111111100000000000000111111",
 "11111000011111110000000000011111110000001111100011111111000000000011111110000000111100001111111000000000000000000000000111100001111111100000000001111111000000011111111111000111111100000000000000111111",
 "11111000011111110000000000000000000000001111100011111111000000000011111110000000111100001111111000000000000000000000000111100001111111100000000001111111000000011111111111000111111100000000000000111111",
 "11111000011111110000000000000000000000001111100011111111000000000011111110000000111100001111111000000000000000000000000111100001111111100000000001111111000000011111111111000111111100000000000000111111",
 "11111000011111110000000000000000000000001111100011111111000000000011111110000000111100001111111000000000000000000000000111100001111111100000000001111111000000011111111111000111111100000000000000011111",
 "11111000011111110000000000000000000000001111100011111111000000000011111110000000111100001111111000000000000000000000000111100001111111100000000001111111000000011111111111000111111100000001111111111111",
 "11111000011111110000000111111111110000001111100011111111111111111111110000000000111100001111111111111111111110000000111111100001111111100000000001111111000000011111111111000111111100000001111111111111",
 "11111000011111110000000111111111110000001111100011111111111111111111110000000000111100001111111111111111111110000000111111100001111111100000000001111111000000011111111111000111111100000001111111111111",
 "11111000011111110000000111111111110000001111100011111111111111111111110000000000111100001111111111111111111110000000111111100001111111000000000001111111000000011111111111000111111100000001111111111111",
 "11111000011111110000000111111111110000001111100011111111111111111111110000000000111100001111111111111111111110000000111111100001111111111111111111111111000000011111111111000111111100000001111111111111",
 "11111000011111110000000000111111110000001111100011111111000000000011111110000000111100001111111000000000000000000000111111100001111111111111111111111111000000011111111111000111111100000001111111111111",
 "11111000011111110000000000011111110000001111100011111111000000000011111110000000111100001111111000000000000000000000111111100001111111111111111111111111000000011111111111000111111100000001111111111111",
 "11111000011111110000000000011111110000001111100011111111000000000011111110000000111100001111111000000000000000000000111111100001111111111111111111111111000000011111111111000111111100000001111111111111",
 "11111000011111110000000000011111110000001111100011111111000000000011111110000000111100001111111000000000000000000000111111100001111111111111111111111111000000011111111111000111111100000001111111111111",
 "11111000011111110000000000011111110000001111100011111111000000000011111110000000111100001111111000000000000000000000111111100001111111100000000001111111000000011111111111000111111100000001111111111111",
 "11111000011111110000000000011111110000001111100011111111000000000011111110000000111100001111111000000000000000000000111111100001111111100000000001111111000000011111111111000111111100000001111111111111",
 "11111000011111110000000000011111110000001111100011111111000000000011111110000000111100001111111000000000000000000000111111100001111111100000000001111111000000011111111111000111111100000001111111111111",
 "11111000011111110000000000011111110000001111100011111111000000000011111110000000111100001111111000000000000000000000111111100001111111100000000001111111000000011111111111000111111100000001111111111111",
 "11111000011111110000000000111111110000001111100011111111000000000011111110000000111100001111111000000000000000000000111111100001111111100000000001111111000000011111111111000111111100000001111111111111",
 "11111000000011111111111111100011110000001111100011111111000000000011111110000000111100001111111111111111111111111000000111100001111111100000000001111111000000011111111111000111111100000001111111111111",
 "11111000000011111111111111100011110000001111100011111111000000000011111110000000111100001111111111111111111111111000000111100001111111100000000001111111000000011111111111000111111100000001111111111111",
 "11111000000011111111111111100011110000001111100011111111000000000011111110000000111100001111111111111111111111111000000111100001111111100000000001111111000000011111111111000111111100000001111111111111",
 "11111000000011111111111111100011110000001111100011111111000000000011111110000000111100001111111111111111111111111000000111100001111111100000000001111111000000011111111111000111111100000001111111111111",
 "11111000000011111111111111100011110000001111100011111111000000000011111110000000111100001111111111111111111111111000000111100000000000000000000000000000000000011111111111000000000000000001111111111111",
 "11111111100000000000000000000000000000001111100000000000000000000000000000000000111100000000000000000000000000000000000111100000000000000000000000000000000000011111111111000000000000000001111111111111",
 "11111111100000000000000000000000000000001111100000000000000000000000000000000000111100000000000000000000000000000000000111100000000000000000000000000000000000011111111111000000000000000001111111111111",
 "11111111100000000000000000000000000000001111100000000000000000000000000000000000111100000000000000000000000000000000000111100000000000000000000000000000000000011111111111000000000000000001111111111111",
 "11111111100000000000000000000000000000001111100000000000000000000000000000000000111100000000000000000000000000000000000111111110000000000000011110000000000000011111111111111000000000000001111111111111",
 "11111111111100000000000000000000000000001111111100000000000000111100000000000000111111110000000000000000000000000000000111111110000000000000011110000000000000011111111111111000000000000001111111111111",
 "11111111111100000000000000000000000000001111111100000000000000111100000000000000111111110000000000000000000000000000000111111110000000000000011110000000000000011111111111111000000000000001111111111111",
 "11111111111100000000000000000000000000001111111100000000000000111100000000000000111111110000000000000000000000000000000111111110000000000000011110000000000000011111111111111000000000000001111111111111",
 "11111111111100000000000000000000000000001111111100000000000000111100000000000000111111110000000000000000000000000000000111111111000000000000011110000000000000011111111111111100000000000001111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");














               
Zero <=                
       ("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
        "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
        "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
        "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
        "111111111111111111111111111111111111000000000000000000111111111111111111111111111111111111",
        "111111111111111111111111111111111110000000000000000000011111111111111111111111111111111111",
        "111111111111111111111111111111111110000000000000000000011111111111111111111111111111111111",
        "111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111",
        "111111111111111111111111111111111000001111111111111000000011111111111111111111111111111111",
        "111111111111111111111111111111111000001111000000011100000001111111111111111111111111111111",
        "111111111111111111111111111111111000111110000000011111000000111111111111111111111111111111",
        "111111111111111111111111111111111000111110000000011111000000111111111111111111111111111111",
        "111111111111111111111111111111111000111110000000011111000000111111111111111111111111111111",
        "111111111111111111111111111111111000111110000001111111000000111111111111111111111111111111",
        "111111111111111111111111111111111000111110000001111111000000111111111111111111111111111111",
        "111111111111111111111111111111111000111110001100011111000000111111111111111111111111111111",
        "111111111111111111111111111111111000111110001100011111000000111111111111111111111111111111",
        "111111111111111111111111111111111000111110000100011111000000111111111111111111111111111111",
        "111111111111111111111111111111111000111111100000011111000000111111111111111111111111111111",
        "111111111111111111111111111111111000111111100000011111000000111111111111111111111111111111",
        "111111111111111111111111111111111000111110000000011111000000111111111111111111111111111111",
        "111111111111111111111111111111111000111110000000011111000000111111111111111111111111111111",
        "111111111111111111111111111111111000111110000000011111000000111111111111111111111111111111",
        "111111111111111111111111111111111000001111111111111100000000111111111111111111111111111111",
        "111111111111111111111111111111111000001111111111111000000000111111111111111111111111111111",
        "111111111111111111111111111111111000001111111111111000000000111111111111111111111111111111",
        "111111111111111111111111111111111110000000000000000000000000111111111111111111111111111111",
        "111111111111111111111111111111111110000000000000000000000000111111111111111111111111111111",
        "111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111",
        "111111111111111111111111111111111111110000000000000000000011111111111111111111111111111111",
        "111111111111111111111111111111111111110000000000000000000011111111111111111111111111111111",
        "111111111111111111111111111111111111111000000000000000000111111111111111111111111111111111",
        "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
        "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111",
        "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");

One <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111110000000000011111111111111111111111111111111111111111", 
 "111111111111111111111111111111111110000000000000000111111111111111111111111111111111111111", 
 "111111111111111111111111111111111110000001111100000111111111111111111111111111111111111111", 
 "111111111111111111111111111111111110000001111100000111111111111111111111111111111111111111", 
 "111111111111111111111111111111111110000011111100000111111111111111111111111111111111111111", 
 "111111111111111111111111111111111110001111111100000111111111111111111111111111111111111111", 
 "111111111111111111111111111111111110001011111100000111111111111111111111111111111111111111", 
 "111111111111111111111111111111111110000001111100000111111111111111111111111111111111111111", 
 "111111111111111111111111111111111110000001111100000111111111111111111111111111111111111111", 
 "111111111111111111111111111111111110000001111100000111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111110001111100000111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111110001111100000111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111110001111100000111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111110001111100000111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111100001111100000111111111111111111111111111111111111111", 
 "111111111111111111111111111111110000000001111100000000111111111111111111111111111111111111", 
 "111111111111111111111111111111110000000001111100000000111111111111111111111111111111111111", 
 "111111111111111111111111111111110000000001111100000000011111111111111111111111111111111111", 
 "111111111111111111111111111111110001111111111111111000000111111111111111111111111111111111", 
 "111111111111111111111111111111110000111111111111111000000111111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111", 
 "111111111111111111111111111111111000000000000000000000000111111111111111111111111111111111", 
 "111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111", 
 "111111111111111111111111111111111110000000000000000000000111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");

Two <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111", 
 "111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111", 
 "111111111111111111111111111111110000001111111111111000000111111111111111111111111111111111", 
 "111111111111111111111111111111110000001111111111111000000111111111111111111111111111111111", 
 "111111111111111111111111111111110000011100000000011000000001111111111111111111111111111111", 
 "111111111111111111111111111111110001111100000000011110000001111111111111111111111111111111", 
 "111111111111111111111111111111110001111100000000011110000001111111111111111111111111111111", 
 "111111111111111111111111111111110001111100000011111110000001111111111111111111111111111111", 
 "111111111111111111111111111111110001111100000011111110000001111111111111111111111111111111", 
 "111111111111111111111111111111110000111100000011111110000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000011111111000000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000011111111000000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000011111000000000001111111111111111111111111111111", 
 "111111111111111111111111111111111110000001111111000000000001111111111111111111111111111111", 
 "111111111111111111111111111111111100000001111111000000000001111111111111111111111111111111", 
 "111111111111111111111111111111110000001111111000000000000011111111111111111111111111111111", 
 "111111111111111111111111111111110000001111111000000000000111111111111111111111111111111111", 
 "111111111111111111111111111111110000001111111000000000000111111111111111111111111111111111", 
 "111111111111111111111111111111110001111111111111111110000001111111111111111111111111111111", 
 "111111111111111111111111111111110001111111111111111110000001111111111111111111111111111111", 
 "111111111111111111111111111111110000010000000000000100000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000000000000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000000000000001111111111111111111111111111111", 
 "111111111111111111111111111111111000000000000000000000000001111111111111111111111111111111", 
 "111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111", 
 "111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");


Three <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111", 
 "111111111111111111111111111111111110000000000000000000111111111111111111111111111111111111", 
 "111111111111111111111111111111111100000000000000000000111111111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111", 
 "111111111111111111111111111111110000001111111111111000000111111111111111111111111111111111", 
 "111111111111111111111111111111110000001110000000111000000001111111111111111111111111111111", 
 "111111111111111111111111111111110001111100000000011110000001111111111111111111111111111111", 
 "111111111111111111111111111111110001111100000000011110000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000011110000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000011110000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000011110000001111111111111111111111111111111", 
 "111111111111111111111111111111111110000000011111111000000001111111111111111111111111111111", 
 "111111111111111111111111111111111110000000011111111000000001111111111111111111111111111111", 
 "111111111111111111111111111111111100000000001111111000000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000011110000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000011110000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000011110000001111111111111111111111111111111", 
 "111111111111111111111111111111110001111100000000011110000001111111111111111111111111111111", 
 "111111111111111111111111111111110001111100000000011110000001111111111111111111111111111111", 
 "111111111111111111111111111111110000001111111111111000000001111111111111111111111111111111", 
 "111111111111111111111111111111110000001111111111111000000001111111111111111111111111111111", 
 "111111111111111111111111111111110000001111111111111000000001111111111111111111111111111111", 
 "111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111", 
 "111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111", 
 "111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111", 
 "111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111", 
 "111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111", 
 "111111111111111111111111111111111111110000000000000000001111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");

Four <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111110000000000011111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111100000000000011111111111111111111111111111111111", 
 "111111111111111111111111111111111111111110000000000000000011111111111111111111111111111111", 
 "111111111111111111111111111111111111111110000001111100000011111111111111111111111111111111", 
 "111111111111111111111111111111111111111110000001111100000011111111111111111111111111111111", 
 "111111111111111111111111111111111111110000001111111100000011111111111111111111111111111111", 
 "111111111111111111111111111111111111110000001111111100000011111111111111111111111111111111", 
 "111111111111111111111111111111111111000000001111111100000011111111111111111111111111111111", 
 "111111111111111111111111111111111111000000111111111100000011111111111111111111111111111111", 
 "111111111111111111111111111111111110000000111111111100000011111111111111111111111111111111", 
 "111111111111111111111111111111111000000111110001111100000011111111111111111111111111111111", 
 "111111111111111111111111111111111000000111110001111100000011111111111111111111111111111111", 
 "111111111111111111111111111111111000000111100001111100000011111111111111111111111111111111", 
 "111111111111111111111111111111111000111110000001111100000011111111111111111111111111111111", 
 "111111111111111111111111111111111000111110000001111100000011111111111111111111111111111111", 
 "111111111111111111111111111111111000111111000011111100000000111111111111111111111111111111", 
 "111111111111111111111111111111111000111111111111111111000000111111111111111111111111111111", 
 "111111111111111111111111111111111000111111111111111111000000111111111111111111111111111111", 
 "111111111111111111111111111111111000000000000001111100000000111111111111111111111111111111", 
 "111111111111111111111111111111111000000000000001111100000000111111111111111111111111111111", 
 "111111111111111111111111111111111000000000000001111100000000111111111111111111111111111111", 
 "111111111111111111111111111111111110000000000000000000000000111111111111111111111111111111", 
 "111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111", 
 "111111111111111111111111111111111111000000000000000000000000111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111100000000000011111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");

Five <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000000000000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000000000000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000000000000001111111111111111111111111111111", 
 "111111111111111111111111111111110001111111111111111110000001111111111111111111111111111111", 
 "111111111111111111111111111111110001111111111111111110000001111111111111111111111111111111", 
 "111111111111111111111111111111110001111100000000000000000001111111111111111111111111111111", 
 "111111111111111111111111111111110001111100000000000000000001111111111111111111111111111111", 
 "111111111111111111111111111111110001111100000000000000000001111111111111111111111111111111", 
 "111111111111111111111111111111110001111111111111111000000001111111111111111111111111111111", 
 "111111111111111111111111111111110001111111111111111000000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000111000000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000011110000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000011110000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000011110000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000011110000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000011110000001111111111111111111111111111111", 
 "111111111111111111111111111111110000111100000000011110000001111111111111111111111111111111", 
 "111111111111111111111111111111110001111100000000011110000001111111111111111111111111111111", 
 "111111111111111111111111111111110000111100000000111110000001111111111111111111111111111111", 
 "111111111111111111111111111111110000001111111111111000000001111111111111111111111111111111", 
 "111111111111111111111111111111110000001111111111111000000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000000000000001111111111111111111111111111111", 
 "111111111111111111111111111111111100000000000000000000000001111111111111111111111111111111", 
 "111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111", 
 "111111111111111111111111111111111110000000000000000000000001111111111111111111111111111111", 
 "111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111", 
 "111111111111111111111111111111111111100000000000000000000111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");

Six <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111100000000000001111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111100000000000001111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111000000000000001111111111111111111111111111111111111111", 
 "111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111", 
 "111111111111111111111111111111111100000011111110000001111111111111111111111111111111111111", 
 "111111111111111111111111111111110000000011100000000001111111111111111111111111111111111111", 
 "111111111111111111111111111111100000011111000000000001111111111111111111111111111111111111", 
 "111111111111111111111111111111100000011111000000000001111111111111111111111111111111111111", 
 "111111111111111111111111111111100000111100000000000001111111111111111111111111111111111111", 
 "111111111111111111111111111111100001111000000000000001111111111111111111111111111111111111", 
 "111111111111111111111111111111100001111100000000000001111111111111111111111111111111111111", 
 "111111111111111111111111111111100011111111111111110000001111111111111111111111111111111111", 
 "111111111111111111111111111111100001111111111111110000001111111111111111111111111111111111", 
 "111111111111111111111111111111100001111100000001110000000011111111111111111111111111111111", 
 "111111111111111111111111111111100001111000000000111110000011111111111111111111111111111111", 
 "111111111111111111111111111111100001111000000000111110000011111111111111111111111111111111", 
 "111111111111111111111111111111100001111000000000111110000011111111111111111111111111111111", 
 "111111111111111111111111111111100001111000000000111110000011111111111111111111111111111111", 
 "111111111111111111111111111111100001111000000000111110000011111111111111111111111111111111", 
 "111111111111111111111111111111100000011111111111110000000011111111111111111111111111111111", 
 "111111111111111111111111111111100000011111111111110000000011111111111111111111111111111111", 
 "111111111111111111111111111111100000011111111111110000000011111111111111111111111111111111", 
 "111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111", 
 "111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111", 
 "111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111", 
 "111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111", 
 "111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111", 
 "111111111111111111111111111111111111110001111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");

Seven <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000000000001111111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000000000000111111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000000000000001111111111111111111111111111111", 
 "111111111111111111111111111111110001111111111111111110000001111111111111111111111111111111", 
 "111111111111111111111111111111110001111111111111111110000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000011111000000001111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000011111000000001111111111111111111111111111111", 
 "111111111111111111111111111111111000000000000011111000000001111111111111111111111111111111", 
 "111111111111111111111111111111111110000000000011111000000001111111111111111111111111111111", 
 "111111111111111111111111111111111110000000000011111000000001111111111111111111111111111111", 
 "111111111111111111111111111111111111111100001111000000000111111111111111111111111111111111", 
 "111111111111111111111111111111111111111100011111000000000111111111111111111111111111111111", 
 "111111111111111111111111111111111111111100011111000000000111111111111111111111111111111111", 
 "111111111111111111111111111111111111100000011111000000000111111111111111111111111111111111", 
 "111111111111111111111111111111111111100000011111000000000111111111111111111111111111111111", 
 "111111111111111111111111111111111111100000011000000000001111111111111111111111111111111111", 
 "111111111111111111111111111111111111100001111000000000111111111111111111111111111111111111", 
 "111111111111111111111111111111111111100001111000000000111111111111111111111111111111111111", 
 "111111111111111111111111111111111111100001111000000000111111111111111111111111111111111111", 
 "111111111111111111111111111111111111100001111000000000111111111111111111111111111111111111", 
 "111111111111111111111111111111111111100000000000000000111111111111111111111111111111111111", 
 "111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111100000000000000111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111110000000000000111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111100000000000111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");

Eight <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111110010000000000001011111111111111111111111111111111111111", 
 "111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111", 
 "111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111", 
 "111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111", 
 "111111111111111111111111111111100000011111111111110000001111111111111111111111111111111111", 
 "111111111111111111111111111111100001111100000000111100000011111111111111111111111111111111", 
 "111111111111111111111111111111100001111000000000111110000011111111111111111111111111111111", 
 "111111111111111111111111111111100001111100000000111110000011111111111111111111111111111111", 
 "111111111111111111111111111111100001111100000000111110000011111111111111111111111111111111", 
 "111111111111111111111111111111100001111111000000111110000011111111111111111111111111111111", 
 "111111111111111111111111111111100001111111000000111110000011111111111111111111111111111111", 
 "111111111111111111111111111111100000011111100001110000000011111111111111111111111111111111", 
 "111111111111111111111111111111100000011111111111110000000011111111111111111111111111111111", 
 "111111111111111111111111111111100000011111111111110000000011111111111111111111111111111111", 
 "111111111111111111111111111111100001111100000111111100000011111111111111111111111111111111", 
 "111111111111111111111111111111100001111000000111111110000011111111111111111111111111111111", 
 "111111111111111111111111111111100001111000000001111110000011111111111111111111111111111111", 
 "111111111111111111111111111111100001111000000000111110000011111111111111111111111111111111", 
 "111111111111111111111111111111100001111000000000111110000011111111111111111111111111111111", 
 "111111111111111111111111111111100000011100000000111000000011111111111111111111111111111111", 
 "111111111111111111111111111111100000011111111111110000000011111111111111111111111111111111", 
 "111111111111111111111111111111100000011111111111110000000011111111111111111111111111111111", 
 "111111111111111111111111111111110000000000000000000000000011111111111111111111111111111111", 
 "111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111", 
 "111111111111111111111111111111111100000000000000000000000011111111111111111111111111111111", 
 "111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111", 
 "111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111", 
 "111111111111111111111111111111111111100000000000000000001111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");

Nine <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111", 
 "111111111111111111111111111111111100000000000000000001111111111111111111111111111111111111", 
 "111111111111111111111111111111111000000000000000000001111111111111111111111111111111111111", 
 "111111111111111111111111111111100000000000000000000000001111111111111111111111111111111111", 
 "111111111111111111111111111111100000011111111111110000001111111111111111111111111111111111", 
 "111111111111111111111111111111100000011100000001110000000011111111111111111111111111111111", 
 "111111111111111111111111111111100011111000000000111100000011111111111111111111111111111111", 
 "111111111111111111111111111111100011111000000000111100000011111111111111111111111111111111", 
 "111111111111111111111111111111100011111000000000111100000011111111111111111111111111111111", 
 "111111111111111111111111111111100011111000000000111100000011111111111111111111111111111111", 
 "111111111111111111111111111111100011111000000000111100000011111111111111111111111111111111", 
 "111111111111111111111111111111100000011111111111111100000011111111111111111111111111111111", 
 "111111111111111111111111111111100000011111111111111100000011111111111111111111111111111111", 
 "111111111111111111111111111111100000011111111111111100000011111111111111111111111111111111", 
 "111111111111111111111111111111111100000000000000111100000011111111111111111111111111111111", 
 "111111111111111111111111111111111100000000000000111100000011111111111111111111111111111111", 
 "111111111111111111111111111111111100000000000001110000000011111111111111111111111111111111", 
 "111111111111111111111111111111111111000000000111110000000011111111111111111111111111111111", 
 "111111111111111111111111111111111111000000000111110000000011111111111111111111111111111111", 
 "111111111111111111111111111111111111000011111110000000000011111111111111111111111111111111", 
 "111111111111111111111111111111111111000011111110000000000011111111111111111111111111111111", 
 "111111111111111111111111111111111111000011111110000000000011111111111111111111111111111111", 
 "111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111", 
 "111111111111111111111111111111111111000000000000000000001111111111111111111111111111111111", 
 "111111111111111111111111111111111111100000000000000000011111111111111111111111111111111111", 
 "111111111111111111111111111111111111111000000000000001111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111100000000000001111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");

Ten <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111110000000000001111111111111111110000000000000000001111111111111111111111", 
 "111111111111111111110000000000001111111111111111100000000000000000000111111111111111111111", 
 "111111111111111111000000000000000011111111111111100000000000000000000111111111111111111111", 
 "111111111111111111000000111100000011111111111110000000000000000000000001111111111111111111", 
 "111111111111111111000000111100000011111111111110000011111111111110000000111111111111111111", 
 "111111111111111111000111111100000011111111111110000011100000001110000000011111111111111111", 
 "111111111111111111000111111100000011111111111110001111100000000111110000001111111111111111", 
 "111111111111111111000001111100000011111111111110001111100000000111110000001111111111111111", 
 "111111111111111111000000111100000011111111111110001111100000000111110000001111111111111111", 
 "111111111111111111000000111100000011111111111110001111100000011111110000001111111111111111", 
 "111111111111111111100000111100000011111111111110001111100000011111110000001111111111111111", 
 "111111111111111111110000111100000011111111111110001111100011000111110000001111111111111111", 
 "111111111111111111110000111100000011111111111110001111100011000111110000001111111111111111", 
 "111111111111111111110000111100000011111111111110001111100010000111110000001111111111111111", 
 "111111111111111111110000111100000011111111111110001111111000000111110000001111111111111111", 
 "111111111111111000000000111100000000011111111110001111111000000111110000001111111111111111", 
 "111111111111111000000000111100000000011111111110001111100000000111110000001111111111111111", 
 "111111111111111000000000111100000000011111111110001111100000000111110000001111111111111111", 
 "111111111111111000000001111110000000000111111110001111100000000111110000001111111111111111", 
 "111111111111111000111111111111111100000011111110000011111111111111000000001111111111111111", 
 "111111111111111000111111111111111100000011111110000011111111111110000000001111111111111111", 
 "111111111111111000000000000000000000000011111110000011111111111110000000001111111111111111", 
 "111111111111111000000000000000000000000011111111100000000000000000000000001111111111111111", 
 "111111111111111000000000000000000000000011111111100000000000000000000000001111111111111111", 
 "111111111111111110000000000000000000000011111111100000000000000000000000001111111111111111", 
 "111111111111111111000000000000000000000011111111111100000000000000000000111111111111111111", 
 "111111111111111111000000000000000000000011111111111100000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");

Eleven       <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111110000000000111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111100000000000111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111100000000000011111111111111111111000000000000111111111111111111111111", 
 "111111111111111111100000000000000000111111111111111111000000000000111111111111111111111111", 
 "111111111111111111100000011111000000111111111111111100000000000000001111111111111111111111", 
 "111111111111111111100000011111000000111111111111111100000011110000001111111111111111111111", 
 "111111111111111111100011111111000000111111111111111100000011110000001111111111111111111111", 
 "111111111111111111100001111111000000111111111111111100000111110000001111111111111111111111", 
 "111111111111111111100000011111000000111111111111111100011111110000001111111111111111111111", 
 "111111111111111111100000011111000000111111111111111100000111110000001111111111111111111111", 
 "111111111111111111100000011111000000111111111111111100000011110000001111111111111111111111", 
 "111111111111111111111100011111000000111111111111111100000011110000001111111111111111111111", 
 "111111111111111111111100011111000000111111111111111100000011110000001111111111111111111111", 
 "111111111111111111111100011111000000111111111111111111000011110000001111111111111111111111", 
 "111111111111111111111100011111000000111111111111111111000011110000001111111111111111111111", 
 "111111111111111111111100011111000000111111111111111111000011110000001111111111111111111111", 
 "111111111111111110000000011111000000000111111111111111000011110000001111111111111111111111", 
 "111111111111111110000000011111000000000111111111111111000011110000001111111111111111111111", 
 "111111111111111110000000011111000000000111111111100000000011110000000001111111111111111111", 
 "111111111111111110000010011111100000000001111111100000000011110000000001111111111111111111", 
 "111111111111111110001111111111111110000000111111100000000011111000000001111111111111111111", 
 "111111111111111110001111111111111110000000111111100011111111111111110000001111111111111111", 
 "111111111111111110000000000000000000000000111111100011111111111111110000001111111111111111", 
 "111111111111111110000000000000000000000000111111100000000000000000000000001111111111111111", 
 "111111111111111110000000000000000000000000111111100000000000000000000000001111111111111111", 
 "111111111111111111100000000000000000000000111111100000000000000000000000001111111111111111", 
 "111111111111111111100000000000000000000000111111110000000000000000000000001111111111111111", 
 "111111111111111111110000000000000000000001111111111100000000000000000000001111111111111111", 
 "111111111111111111111111111111111111111111111111111100000000000000000000001111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Twelve       <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111100000000000111111111111111110000000000000000000111111111111111111111", 
 "111111111111111111111100000000000111111111111111100000000000000000000111111111111111111111", 
 "111111111111111111110000000000000001111111111110000000000000000000000001111111111111111111", 
 "111111111111111111100000011111000000111111111110000001111111111110000000111111111111111111", 
 "111111111111111111100000011111000000111111111110000001111111111110000000111111111111111111", 
 "111111111111111111100000011111000000111111111110000011100000000111000000001111111111111111", 
 "111111111111111111100011111111000000111111111110001111100000000011110000001111111111111111", 
 "111111111111111111100001111111000000111111111110001111100000000111110000001111111111111111", 
 "111111111111111111100000011111000000111111111110001111100000011111110000001111111111111111", 
 "111111111111111111100000011111000000111111111110001111100000011111110000001111111111111111", 
 "111111111111111111110000011111000000111111111110000111100000011111110000001111111111111111", 
 "111111111111111111111100011111000000111111111110000000000011111111000000001111111111111111", 
 "111111111111111111111100011111000000111111111110000000000011111110000000001111111111111111", 
 "111111111111111111111100011111000000111111111110000000000011111000000000001111111111111111", 
 "111111111111111111111100011111000000111111111111100000011111111000000000001111111111111111", 
 "111111111111111111111100011111000000111111111111100000011111110000000000001111111111111111", 
 "111111111111111110000000011111000000000111111110000001111111000000000000111111111111111111", 
 "111111111111111110000000011111000000000111111110000001111111000000000000111111111111111111", 
 "111111111111111110000000011111000000000111111110000001111111000000000000111111111111111111", 
 "111111111111111110001111111111111110000000111110001111111111111111110000001111111111111111", 
 "111111111111111110001111111111111110000000111110001111111111111111110000001111111111111111", 
 "111111111111111110000010000000000000000000111110000010000000000001000000001111111111111111", 
 "111111111111111110000000000000000000000000111110000000000000000000000000001111111111111111", 
 "111111111111111110000000000000000000000000111110000000000000000000000000001111111111111111", 
 "111111111111111110000000000000000000000000111110000000000000000000000000001111111111111111", 
 "111111111111111111100000000000000000000000111111100000000000000000000000001111111111111111", 
 "111111111111111111100000000000000000000000111111110000000000000000000000001111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Thirteen     <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111000000000011111111111111111000000000000000000011111111111111111111", 
 "111111111111111111111110000000000011111111111111110000000000000000000011111111111111111111", 
 "111111111111111111111110000000000001111111111111110000000000000000000011111111111111111111", 
 "111111111111111111110000000000000000011111111111000000000000000000000000011111111111111111", 
 "111111111111111111110000001111100000011111111111000000111111111111000000011111111111111111", 
 "111111111111111111110000001111100000011111111111000001110000000011100000000111111111111111", 
 "111111111111111111110001111111100000011111111111000111110000000001111000000111111111111111", 
 "111111111111111111110000111111100000011111111111000011110000000001111000000111111111111111", 
 "111111111111111111110000001111100000011111111111000000000000000001111000000111111111111111", 
 "111111111111111111110000001111100000011111111111000000000000000001111000000111111111111111", 
 "111111111111111111110000001111100000011111111111000000000000000001111000000111111111111111", 
 "111111111111111111111110001111100000011111111111111000000001111111100000000111111111111111", 
 "111111111111111111111110001111100000011111111111110000000001111111000000000111111111111111", 
 "111111111111111111111110001111100000011111111111110000000000111111100000000111111111111111", 
 "111111111111111111111110001111100000011111111111000000000000000001111000000111111111111111", 
 "111111111111111111111110001111100000011111111111000000000000000001111000000111111111111111", 
 "111111111111111111000000001111100000000011111111000000000000000001111000000111111111111111", 
 "111111111111111111000000001111100000000011111111000111110000000001111000000111111111111111", 
 "111111111111111111000000001111100000000011111111000111110000000001111000000111111111111111", 
 "111111111111111111000011111111111111000000111111000001111111111111100000000111111111111111", 
 "111111111111111111000111111111111111000000011111000000111111111111100000000111111111111111", 
 "111111111111111111000111111111111111000000011111000000111111111111000000000111111111111111", 
 "111111111111111111000000000000000000000000011111110000000000000000000000000111111111111111", 
 "111111111111111111000000000000000000000000011111110000000000000000000000000111111111111111", 
 "111111111111111111000000000000000000000000011111111000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000011111111110000000000000000000011111111111111111", 
 "111111111111111111110000000000000000000000011111111110000000000000000000011111111111111111", 
 "111111111111111111111000000000000000000000111111111111000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Fourteen     <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111100000000000111111111111111111111111100000000000111111111111111111111", 
 "111111111111111111111100000000000111111111111111111111111100000000000111111111111111111111", 
 "111111111111111111111100000000000011111111111111111111111000000000000111111111111111111111", 
 "111111111111111111100000000000000000111111111111111111100000000000000000111111111111111111", 
 "111111111111111111100000011111000000111111111111111111100000011110000000111111111111111111", 
 "111111111111111111100000011111000000111111111111111111100000011110000000111111111111111111", 
 "111111111111111111100011111111000000111111111111111100000011111110000000111111111111111111", 
 "111111111111111111100001111111000000111111111111111100000011111110000000111111111111111111", 
 "111111111111111111100000011111000000111111111111110000000011111110000000111111111111111111", 
 "111111111111111111100000011111000000111111111111100000011111111110000000111111111111111111", 
 "111111111111111111100000011111000000111111111111100000011111111111000000111111111111111111", 
 "111111111111111111111100011111000000111111111110000001111100011111000000111111111111111111", 
 "111111111111111111111100011111000000111111111110000001111100011111000000111111111111111111", 
 "111111111111111111111100011111000000111111111110000001111000011110000000111111111111111111", 
 "111111111111111111111100011111000000111111111110001111100000011110000000111111111111111111", 
 "111111111111111111111100011111000000111111111110001111100000011110000000111111111111111111", 
 "111111111111111110000000011111000000000111111110001111100000111111000000001111111111111111", 
 "111111111111111110000000011111000000000111111110001111111111111111110000001111111111111111", 
 "111111111111111110000000011111000000000111111110001111111111111111110000001111111111111111", 
 "111111111111111110000111111111111110000001111110000000000000011111000000001111111111111111", 
 "111111111111111110001111111111111110000000111110000000000000011110000000001111111111111111", 
 "111111111111111110001111111111111110000000111110000000000000011110000000001111111111111111", 
 "111111111111111110000000000000000000000000111111100000000000000000000000001111111111111111", 
 "111111111111111110000000000000000000000000111111100000000000000000000000001111111111111111", 
 "111111111111111110000000000000000000000000111111110000000000000000000000001111111111111111", 
 "111111111111111111100000000000000000000000111111111111111111000000000000111111111111111111", 
 "111111111111111111100000000000000000000000111111111111111111000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Fifteen      <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111100000000000111111111111110000000000000000000000000001111111111111111", 
 "111111111111111111111100000000000111111111111110000000000000000000000000001111111111111111", 
 "111111111111111111110000000000000001111111111110000000000000000000000000001111111111111111", 
 "111111111111111111100000011111000000111111111110000111111111111111110000001111111111111111", 
 "111111111111111111100000011111000000111111111110001111111111111111110000001111111111111111", 
 "111111111111111111100000011111000000111111111110001111100000000000000000001111111111111111", 
 "111111111111111111100011111111000000111111111110001111100000000000000000001111111111111111", 
 "111111111111111111100000011111000000111111111110001111100000000000000000001111111111111111", 
 "111111111111111111100000011111000000111111111110001111111111111110000000001111111111111111", 
 "111111111111111111100000011111000000111111111110001111111111111110000000001111111111111111", 
 "111111111111111111110000011111000000111111111110000000000000000111000000001111111111111111", 
 "111111111111111111111100011111000000111111111110000000000000000011110000001111111111111111", 
 "111111111111111111111100011111000000111111111110000000000000000011110000001111111111111111", 
 "111111111111111111111100011111000000111111111110000000000000000011110000001111111111111111", 
 "111111111111111111111100011111000000111111111110000000000000000011110000001111111111111111", 
 "111111111111111111111100011111000000111111111110000000000000000011110000001111111111111111", 
 "111111111111111110000000011111000000000111111110000111100000000011110000001111111111111111", 
 "111111111111111110000000011111000000000111111110001111100000000011110000001111111111111111", 
 "111111111111111110000000011111000000000111111110000111100000000111110000001111111111111111", 
 "111111111111111110001111111111111110000000111110000001111111111111000000001111111111111111", 
 "111111111111111110001111111111111110000000111110000001111111111110000000001111111111111111", 
 "111111111111111110000000000000000000000000111110000000000000000000000000001111111111111111", 
 "111111111111111110000000000000000000000000111111100000000000000000000000001111111111111111", 
 "111111111111111110000000000000000000000000111111100000000000000000000000001111111111111111", 
 "111111111111111111000000000000000000000000111111111000000000000000000000011111111111111111", 
 "111111111111111111100000000000000000000000111111111100000000000000000000111111111111111111", 
 "111111111111111111100000000000000000000000111111111100000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Sixteen      <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111100000000000111111111111111111000000000000011111111111111111111111111", 
 "111111111111111111111100000000000111111111111111110000000000000011111111111111111111111111", 
 "111111111111111111100000000000000001111111111111110000000000000001111111111111111111111111", 
 "111111111111111111100000011111000001111111111111000000000000000000011111111111111111111111", 
 "111111111111111111100000011111000001111111111111000000111111100000011111111111111111111111", 
 "111111111111111111100011111111000001111111111100000000110000000000011111111111111111111111", 
 "111111111111111111100011111111000001111111111000000111110000000000011111111111111111111111", 
 "111111111111111111100000011111000001111111111000000111110000000000011111111111111111111111", 
 "111111111111111111100000011111000001111111111000001110000000000000011111111111111111111111", 
 "111111111111111111100000011111000001111111111000011110000000000000011111111111111111111111", 
 "111111111111111111111100011111000001111111111000011110000000000000011111111111111111111111", 
 "111111111111111111111100011111000001111111111000111111111111111100000011111111111111111111", 
 "111111111111111111111100011111000001111111111000011111111111111100000011111111111111111111", 
 "111111111111111111111100011111000001111111111000011111000000011100000001111111111111111111", 
 "111111111111111111111100011111000001111111111000011110000000001111100000111111111111111111", 
 "111111111111111110000000011111000000001111111000011110000000001111100000111111111111111111", 
 "111111111111111100000000011111000000000111111000011110000000001111100000111111111111111111", 
 "111111111111111100000000011111000000000111111000011110000000001111100000111111111111111111", 
 "111111111111111110001111111111111110000001111000011110000000001111100000111111111111111111", 
 "111111111111111100001111111111111110000001111000000111111111111100000000111111111111111111", 
 "111111111111111100001111111111111110000001111000000111111111111100000000111111111111111111", 
 "111111111111111100000000000000000000000001111000000111111111111100000000111111111111111111", 
 "111111111111111100000000000000000000000001111111000000000000000000000000111111111111111111", 
 "111111111111111110000000000000000000000001111111000000000000000000000000111111111111111111", 
 "111111111111111111100000000000000000000001111111000000000000000000000000111111111111111111", 
 "111111111111111111100000000000000000000001111111110000000000000000000011111111111111111111", 
 "111111111111111111110000000000000000000001111111110000000000000000000011111111111111111111", 
 "111111111111111111111111111111111111111111111111111000011111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Seventeen    <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111110000000000011111111111100000000000000000000000011111111111111111111", 
 "111111111111111111111110000000000011111111111100000000000000000000000001111111111111111111", 
 "111111111111111111110000000000000000111111111100000000000000000000000001111111111111111111", 
 "111111111111111111110000001111000000111111111100000000000000000000000000011111111111111111", 
 "111111111111111111110000001111000000111111111100011111111111111111100000011111111111111111", 
 "111111111111111111110001111111000000111111111100001111111111111111100000011111111111111111", 
 "111111111111111111110001111111000000111111111100000000000000111100000000011111111111111111", 
 "111111111111111111110000001111000000111111111100000000000000111100000000011111111111111111", 
 "111111111111111111110000001111000000111111111100000000000000111100000000011111111111111111", 
 "111111111111111111110000001111000000111111111111000000000000111100000000011111111111111111", 
 "111111111111111111111000001111100000111111111111100000000000111100000000011111111111111111", 
 "111111111111111111111110001111000000111111111111111111000011110000000001111111111111111111", 
 "111111111111111111111110001111000000111111111111111111000111110000000001111111111111111111", 
 "111111111111111111111110001111000000111111111111111111000111110000000001111111111111111111", 
 "111111111111111111111110001111000000111111111111111000000111110000000001111111111111111111", 
 "111111111111111111000000001111000000000111111111111000000111110000000001111111111111111111", 
 "111111111111111110000000001111000000000111111111111000000110000000000011111111111111111111", 
 "111111111111111110000000001111000000000111111111111000111110000000001111111111111111111111", 
 "111111111111111110000000001111100000000001111111111000111110000000001111111111111111111111", 
 "111111111111111110000111111111111111000000111111111000111110000000001111111111111111111111", 
 "111111111111111110000111111111111111000000111111111000111110000000001111111111111111111111", 
 "111111111111111110000000000000000000000000111111111000000000000000001111111111111111111111", 
 "111111111111111110000000000000000000000000111111111000000000000001111111111111111111111111", 
 "111111111111111110000000000000000000000000111111111000000000000001111111111111111111111111", 
 "111111111111111111110000000000000000000000111111111100000000000001111111111111111111111111", 
 "111111111111111111110000000000000000000000111111111111000000000001111111111111111111111111", 
 "111111111111111111110000000000000000000000111111111111000000000001111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Eighteen     <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111000000000001111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111000000000001111111111111110100000000000001001111111111111111111111", 
 "111111111111111111111100000000000000011111111111100000000000000000001111111111111111111111", 
 "111111111111111111111000000111100000011111111111100000000000000000001111111111111111111111", 
 "111111111111111111111000000111100000011111111100000000000000000000000001111111111111111111", 
 "111111111111111111111000000111100000011111111100000011111111111110000001111111111111111111", 
 "111111111111111111111000111111100000011111111100001111000000000111110000011111111111111111", 
 "111111111111111111111000111111100000011111111100001111000000000111110000011111111111111111", 
 "111111111111111111111000000111100000011111111100001111000000000111110000011111111111111111", 
 "111111111111111111111000000111100000011111111100001111100000000111110000011111111111111111", 
 "111111111111111111111000000111100000011111111100001111111000000111110000011111111111111111", 
 "111111111111111111111111000111110000011111111100001111111000000111110000011111111111111111", 
 "111111111111111111111111000111100000011111111100000011111100001110000000011111111111111111", 
 "111111111111111111111111000111100000011111111100000011111111111110000000011111111111111111", 
 "111111111111111111111111000111100000011111111100000011111111111110000000011111111111111111", 
 "111111111111111111111110000111100000011111111100001111000000111111100000011111111111111111", 
 "111111111111111111000000000111100000000011111100001111000000111111110000011111111111111111", 
 "111111111111111111000000000111100000000011111100001111000000001111110000011111111111111111", 
 "111111111111111111000000000111100000000011111100001111000000000111110000011111111111111111", 
 "111111111111111111000111111111111111100000011100001111000000000111110000011111111111111111", 
 "111111111111111111000011111111111111100000011100000111100000001110000000011111111111111111", 
 "111111111111111111000011111111111111100000011100000011111111111110000000011111111111111111", 
 "111111111111111111000000000000000000000000011100000011111111111110000000011111111111111111", 
 "111111111111111111000000000000000000000000011100000000000000000000000000011111111111111111", 
 "111111111111111111100000000000000000000000011111100000000000000000000000011111111111111111", 
 "111111111111111111111000000000000000000000011111100000000000000000000000011111111111111111", 
 "111111111111111111111000000000000000000000011111111000000000000000000001111111111111111111", 
 "111111111111111111111111111111111111111111111111111000000000000000000001111111111111111111", 
 "111111111111111111111111111111111111111111111111111100000000000000000001111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Nineteen     <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111000000000111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111110000000000011111111111111110000000000000000000111111111111111111111", 
 "111111111111111111111110000000000011111111111111100000000000000000000111111111111111111111", 
 "111111111111111111110000000000000000111111111111100000000000000000000111111111111111111111", 
 "111111111111111111110000001111100000111111111110000000000000000000000000111111111111111111", 
 "111111111111111111110000001111100000111111111110000001111111111110000000111111111111111111", 
 "111111111111111111110001111111100000111111111110000011100000000111000000001111111111111111", 
 "111111111111111111110001111111100000111111111110001111100000000011110000001111111111111111", 
 "111111111111111111110000001111100000111111111110001111100000000011110000001111111111111111", 
 "111111111111111111110000001111100000111111111110001111100000000011110000001111111111111111", 
 "111111111111111111110000001111100000111111111110001111100000000011110000001111111111111111", 
 "111111111111111111111110001111100000111111111110001111100000000111110000001111111111111111", 
 "111111111111111111111110001111100000111111111110000001111111111111110000001111111111111111", 
 "111111111111111111111110001111100000111111111110000001111111111111110000001111111111111111", 
 "111111111111111111111110001111100000111111111110000001111111111111110000001111111111111111", 
 "111111111111111111111110001111100000111111111111100000000000000011110000001111111111111111", 
 "111111111111111111000000001111100000000111111111100000000000000011110000001111111111111111", 
 "111111111111111110000000001111100000000011111111110000000000000111000000001111111111111111", 
 "111111111111111110000000001111100000000011111111111100000000011110000000001111111111111111", 
 "111111111111111111000001001111110000000000111111111100000000011110000000001111111111111111", 
 "111111111111111110000111111111111111000000111111111100001111111000000000001111111111111111", 
 "111111111111111110000111111111111111000000111111111100011111111000000000001111111111111111", 
 "111111111111111110000000000000000000000000111111111100011111111000000000001111111111111111", 
 "111111111111111110000000000000000000000000111111111100000000000000000000111111111111111111", 
 "111111111111111111000000000000000000000000111111111100000000000000000000111111111111111111", 
 "111111111111111111110000000000000000000000111111111110000000000000000001111111111111111111", 
 "111111111111111111110000000000000000000000111111111111100000000000000111111111111111111111", 
 "111111111111111111110000000000000000000000111111111111100000000000000111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Twenty       <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111110000000000000000000011111111111111111111111111111111111111111111111111111", 
 "111111111111111110000000000000000000011111111111111000000000000000000111111111111111111111", 
 "111111111111111000000000000000000000000111111111111000000000000000000011111111111111111111", 
 "111111111111111000000111111111111000000111111111110000000000000000000001111111111111111111", 
 "111111111111111000001111111111111000000011111111000000000000000000000000011111111111111111", 
 "111111111111111000001110000000011100000000111111000000111111111111100000011111111111111111", 
 "111111111111111000111110000000011111000000111111000000111000000011100000000111111111111111", 
 "111111111111111000111110000000011111000000111111000111110000000001111000000111111111111111", 
 "111111111111111000111110000001111111000000111111000111110000000001111000000111111111111111", 
 "111111111111111000111110000001111111000000111111000111110000000011111000000111111111111111", 
 "111111111111111000000000000011111100000000111111000111110000001111111000000111111111111111", 
 "111111111111111000000000001111111000000000111111000111110000001111111000000111111111111111", 
 "111111111111111000000000001111111000000000111111000111110001100001111100000111111111111111", 
 "111111111111111000000000001111100000000000111111000111110001100001111000000111111111111111", 
 "111111111111111110000001111111100000000000111111000111110000100001111000000111111111111111", 
 "111111111111111100000001111111000000000000111111000111111100000001111000000111111111111111", 
 "111111111111111000000111111100000000000011111111000111111110000001111000000111111111111111", 
 "111111111111111000001111111100000000000011111111000111110000000001111000000111111111111111", 
 "111111111111111000001111111100000000000001111111000111110000000001111000000111111111111111", 
 "111111111111111000111111111111111111000000111111000111110000000001111000000111111111111111", 
 "111111111111111000111111111111111111000000111111000000111111111111100000000111111111111111", 
 "111111111111111000000000000000000000000000111111000000111111111111100000000111111111111111", 
 "111111111111111000000000000000000000000000111111000000111111111111100000000111111111111111", 
 "111111111111111000000000000000000000000000111111110000000000000000000000000111111111111111", 
 "111111111111111000000000000000000000000000111111111000000000000000000000000111111111111111", 
 "111111111111111110000000000000000000000000111111111000000000000000000000000111111111111111", 
 "111111111111111110000000000000000000000000111111111110000000000000000000011111111111111111", 
 "111111111111111111111111111111111111111111111111111110000000000000000000011111111111111111", 
 "111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Twenty_One   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111000000000000000000011111111111111111111111111111111111111111111111111111", 
 "111111111111111111000000000000000000001111111111111111110000000000011111111111111111111111", 
 "111111111111111110000000000000000000001111111111111111110000000000011111111111111111111111", 
 "111111111111111100000011111111111100000011111111111111000000000000000111111111111111111111", 
 "111111111111111100000111111111111100000001111111111110000001111100000011111111111111111111", 
 "111111111111111100000111000000001100000000111111111110000001111100000011111111111111111111", 
 "111111111111111100011111000000001111100000011111111110000001111100000011111111111111111111", 
 "111111111111111100011111000000001111100000011111111110001111111100000011111111111111111111", 
 "111111111111111100011111000000111111100000011111111110000011111100000011111111111111111111", 
 "111111111111111100011111000000111111100000011111111110000001111100000011111111111111111111", 
 "111111111111111100011111000001111111100000011111111110000001111100000011111111111111111111", 
 "111111111111111100000000000111111100000000011111111111000001111100000011111111111111111111", 
 "111111111111111100000000000111111100000000011111111111110001111100000011111111111111111111", 
 "111111111111111100000000000111111100000000011111111111110001111100000011111111111111111111", 
 "111111111111111111000000111111110000000000011111111111110001111100000011111111111111111111", 
 "111111111111111111000000111111100000000000011111111111110001111100000011111111111111111111", 
 "111111111111111100000000111110000000000000111111111111110001111100000011111111111111111111", 
 "111111111111111100000111111110000000000001111111111000000001111100000000111111111111111111", 
 "111111111111111100000111111110000000000001111111111000000001111100000000111111111111111111", 
 "111111111111111100011111111111111111100000011111111000000001111100000000011111111111111111", 
 "111111111111111100011111111111111111100000011111111000111111111111111000000111111111111111", 
 "111111111111111100011111111111111111100000011111111000111111111111111000000111111111111111", 
 "111111111111111100000000000000000000000000011111111000000000000000000000000111111111111111", 
 "111111111111111100000000000000000000000000011111111000000000000000000000000111111111111111", 
 "111111111111111100000000000000000000000000011111111000000000000000000000000111111111111111", 
 "111111111111111111000000000000000000000000011111111000000000000000000000000111111111111111", 
 "111111111111111111000000000000000000000000011111111110000000000000000000000111111111111111", 
 "111111111111111111111111111111111111111111111111111110000000000000000000000111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Twenty_Two   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111110000000000000000000111111111111110000000000000000000111111111111111111111", 
 "111111111111111110000000000000000000011111111111110000000000000000000111111111111111111111", 
 "111111111111111000000000000000000000000111111111000000000000000000000000111111111111111111", 
 "111111111111111000000111111111111000000111111110000001111111111111000000111111111111111111", 
 "111111111111111000001111111111111000000011111110000001111111111111000000111111111111111111", 
 "111111111111111000001110000000011100000000111110000001100000000011100000001111111111111111", 
 "111111111111111000111110000000011111000000111110000111100000000011111000001111111111111111", 
 "111111111111111000111110000000011111000000111110000111100000000011111000001111111111111111", 
 "111111111111111000111110000001111111000000111110000111100000011111111000001111111111111111", 
 "111111111111111000111110000001111111000000111110000111100000011111111000001111111111111111", 
 "111111111111111000111100000011111111000000111110000111100000011111110000001111111111111111", 
 "111111111111111000000000001111111000000000111110000000000001111111000000001111111111111111", 
 "111111111111111000000000001111111000000000111110000000000001111111000000001111111111111111", 
 "111111111111111000000000001111100000000000111110000000000011111100000000001111111111111111", 
 "111111111111111110000001111111100000000000111111110000001111111000000000001111111111111111", 
 "111111111111111110000001111111000000000000111111110000001111111000000000001111111111111111", 
 "111111111111111000000111111100000000000011111110000001111111100000000000011111111111111111", 
 "111111111111111000001111111100000000000011111110000001111111100000000000111111111111111111", 
 "111111111111111000001111111100000000000011111110000001111111100000000000111111111111111111", 
 "111111111111111000111111111111111111000000111110000111111111111111111000001111111111111111", 
 "111111111111111000111111111111111111000000111110000111111111111111111000001111111111111111", 
 "111111111111111000001000000000000100000000111110000001000000000000100000001111111111111111", 
 "111111111111111000000000000000000000000000111110000000000000000000000000001111111111111111", 
 "111111111111111000000000000000000000000000111110000000000000000000000000001111111111111111", 
 "111111111111111000000000000000000000000000111111000000000000000000000000001111111111111111", 
 "111111111111111110000000000000000000000000111111110000000000000000000000001111111111111111", 
 "111111111111111110000000000000000000000000111111110000000000000000000000001111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Twenty_Three <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111000000000000000000001111111111111000000000000000000011111111111111111111", 
 "111111111111111111000000000000000000001111111111111000000000000000000011111111111111111111", 
 "111111111111111100000000000000000000000011111111111000000000000000000001111111111111111111", 
 "111111111111111100000111111111111100000001111111000000000000000000000000011111111111111111", 
 "111111111111111100000111111111111100000001111111000000111111111111100000011111111111111111", 
 "111111111111111100011111000000001111100000011111000000111000000011100000000111111111111111", 
 "111111111111111100011111000000001111100000011111000011110000000001111100000111111111111111", 
 "111111111111111100011111000000001111100000011111000011110000000001111100000111111111111111", 
 "111111111111111100011111000000111111100000011111000000000000000001111100000111111111111111", 
 "111111111111111100011111000000111111100000011111000000000000000001111100000111111111111111", 
 "111111111111111100000000000111111110000000011111000000000000000001111100000111111111111111", 
 "111111111111111100000000000111111100000000011111111000000000111111100000000111111111111111", 
 "111111111111111100000000000111111100000000011111111000000000111111100000000111111111111111", 
 "111111111111111111000000011111110000000000011111111000000000111111100000000111111111111111", 
 "111111111111111111000000111111110000000000011111000000000000000001111100000111111111111111", 
 "111111111111111100000000111110000000000000011111000000000000000001111100000111111111111111", 
 "111111111111111100000011111110000000000001111111000000000000000001111100000111111111111111", 
 "111111111111111100000111111110000000000001111111000011110000000001111100000111111111111111", 
 "111111111111111100000111111111000000000000011111000011110000000001111100000111111111111111", 
 "111111111111111100011111111111111111100000011111000000111111111111100000000111111111111111", 
 "111111111111111100011111111111111111100000011111000000111111111111100000000111111111111111", 
 "111111111111111100000000000000000000000000011111000000111111111111100000000111111111111111", 
 "111111111111111100000000000000000000000000011111111000000000000000000000000111111111111111", 
 "111111111111111100000000000000000000000000011111111000000000000000000000000111111111111111", 
 "111111111111111111000000000000000000000000011111111000000000000000000000000111111111111111", 
 "111111111111111111000000000000000000000000011111111111000000000000000000011111111111111111", 
 "111111111111111111100000000000000000000000011111111111000000000000000000011111111111111111", 
 "111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");


Twenty_Four  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111100000000000000000011111111111111111111110000000000011111111111111111111", 
 "111111111111111111000000000000000000001111111111111111111110000000000011111111111111111111", 
 "111111111111111111000000000000000000001111111111111111111110000000000001111111111111111111", 
 "111111111111111100000000000000000000000011111111111111110000000000000000011111111111111111", 
 "111111111111111100000111111111111100000001111111111111110000001111100000011111111111111111", 
 "111111111111111100000111111111111100000001111111111111110000001111100000011111111111111111", 
 "111111111111111100011111000000001111100000011111111111000000111111100000011111111111111111", 
 "111111111111111100011111000000001111100000011111111111000000111111100000011111111111111111", 
 "111111111111111100011111000000001111100000011111111000000001111111100000011111111111111111", 
 "111111111111111100011111000000111111100000011111111000000111111111100000011111111111111111", 
 "111111111111111100011111000001111111100000011111111000000111111111100000011111111111111111", 
 "111111111111111100000000000111111100000000011111000000111110001111100000011111111111111111", 
 "111111111111111100000000000111111100000000011111000000111110001111100000011111111111111111", 
 "111111111111111100000000000111111100000000011111000000111110001111100000011111111111111111", 
 "111111111111111111000000111111110000000000011111000011110000001111100000011111111111111111", 
 "111111111111111111000000111111110000000000011111000011110000001111100000011111111111111111", 
 "111111111111111100000000111110000000000000011111000011111000001111100000000111111111111111", 
 "111111111111111100000111111110000000000001111111000011111111111111111100000111111111111111", 
 "111111111111111100000111111110000000000001111111000011111111111111111100000111111111111111", 
 "111111111111111100011111111111111111100000011111000000000000001111100000000111111111111111", 
 "111111111111111100011111111111111111100000011111000000000000001111100000000111111111111111", 
 "111111111111111100011111111111111111100000011111000000000000001111100000000111111111111111", 
 "111111111111111100000000000000000000000000011111110000000000000000000000000111111111111111", 
 "111111111111111100000000000000000000000000011111111000000000000000000000000111111111111111", 
 "111111111111111100000000000000000000000000011111111000000000000000000000000111111111111111", 
 "111111111111111111000000000000000000000000011111111111111111110000000000011111111111111111", 
 "111111111111111111000000000000000000000000011111111111111111110000000000011111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");


Twenty_Five  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111000000000000000000001111111111000000000000000000000000000111111111111111", 
 "111111111111111111000000000000000000001111111111000000000000000000000000000111111111111111", 
 "111111111111111100000000000000000000000011111111000000000000000000000000000111111111111111", 
 "111111111111111100000011111111111100000011111111000011111111111111111100000111111111111111", 
 "111111111111111100000111111111111100000001111111000011111111111111111100000111111111111111", 
 "111111111111111100000111000000001110000000011111000011111000000000000000000111111111111111", 
 "111111111111111100011111000000001111100000011111000011110000000000000000000111111111111111", 
 "111111111111111100011111000000001111100000011111000011110000000000000000000111111111111111", 
 "111111111111111100011111000000111111100000011111000011111111111111100000000111111111111111", 
 "111111111111111100011111000000111111100000011111000011111111111111100000000111111111111111", 
 "111111111111111100000000000001111110000000011111000000000000000011100000000111111111111111", 
 "111111111111111100000000000111111100000000011111000000000000000001111100000111111111111111", 
 "111111111111111100000000000111111100000000011111000000000000000001111100000111111111111111", 
 "111111111111111100000000000111110000000000011111000000000000000001111100000111111111111111", 
 "111111111111111111000000111111110000000000011111000000000000000001111100000111111111111111", 
 "111111111111111111000000111111100000000000011111000000000000000001111100000111111111111111", 
 "111111111111111100000011111110000000000001111111000011110000000001111100000111111111111111", 
 "111111111111111100000111111110000000000001111111000011110000000001111100000111111111111111", 
 "111111111111111100000111111110000000000001111111000011111000000001111000000111111111111111", 
 "111111111111111100011111111111111111100000011111000000111111111111100000000111111111111111", 
 "111111111111111100011111111111111111100000011111000000111111111111100000000111111111111111", 
 "111111111111111100000000000000000000000000011111000000000000000000000000000111111111111111", 
 "111111111111111100000000000000000000000000011111111000000000000000000000000111111111111111", 
 "111111111111111100000000000000000000000000011111111000000000000000000000000111111111111111", 
 "111111111111111100000000000000000000000000011111111100000000000000000000000111111111111111", 
 "111111111111111111000000000000000000000000011111111111000000000000000000011111111111111111", 
 "111111111111111111000000000000000000000000011111111111000000000000000000011111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");


Twenty_Six   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111100000000000000000000111111111111111000000000000011111111111111111111111", 
 "111111111111111111100000000000000000000111111111111111000000000000001111111111111111111111", 
 "111111111111111110000000000000000000000001111111111110000000000000001111111111111111111111", 
 "111111111111111110000011111111111110000000111111111000000000000000000001111111111111111111", 
 "111111111111111110000011111111111110000000111111111000000111111100000001111111111111111111", 
 "111111111111111110001111100000000111110000001111100000000111000000000001111111111111111111", 
 "111111111111111110001111100000000111110000001111000000111110000000000001111111111111111111", 
 "111111111111111110001111100000000111110000001111000000111110000000000001111111111111111111", 
 "111111111111111110001111100000011111110000001111000001111000000000000001111111111111111111", 
 "111111111111111110001111100000011111110000001111000011111000000000000001111111111111111111", 
 "111111111111111110000000000011111111000000001111000011111000000000000001111111111111111111", 
 "111111111111111110000000000011111110000000001111100011111111111111100000011111111111111111", 
 "111111111111111110000000000011111110000000001111000011111111111111100000011111111111111111", 
 "111111111111111111000000001111111000000000001111000011111100000011100000000111111111111111", 
 "111111111111111111100000011111111000000000001111000011111000000001111100000011111111111111", 
 "111111111111111110000000011111000000000000001111000011111000000001111100000011111111111111", 
 "111111111111111110000001111111000000000000111111000011111000000001111100000011111111111111", 
 "111111111111111110000011111111000000000000111111000011111000000001111100000011111111111111", 
 "111111111111111110001111111111111111110000001111000011111000000001111100000011111111111111", 
 "111111111111111110001111111111111111110000001111100000111111111111100000000011111111111111", 
 "111111111111111110001111111111111111110000001111000000111111111111100000000011111111111111", 
 "111111111111111110000000000000000000000000001111000000111111111111100000000011111111111111", 
 "111111111111111110000000000000000000000000001111111000000000000000000000000011111111111111", 
 "111111111111111110000000000000000000000000001111111000000000000000000000000011111111111111", 
 "111111111111111111100000000000000000000000001111111100000000000000000000000011111111111111", 
 "111111111111111111100000000000000000000000001111111111000000000000000000011111111111111111", 
 "111111111111111111110000000000000000000000001111111111000000000000000000011111111111111111", 
 "111111111111111111111111111111111111111111111111111111100011111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");


Twenty_Seven <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111001000000000000100111111111111111111111111111111111111111111111111111111", 
 "111111111111111110000000000000000000011111111110000000000000000000000000111111111111111111", 
 "111111111111111110000000000000000000011111111110000000000000000000000000111111111111111111", 
 "111111111111111000000000000000000000000111111110000000000000000000000000111111111111111111", 
 "111111111111111000001111111111111000000011111110000000000000000000000000001111111111111111", 
 "111111111111111000001111111111111000000011111110000111111111111111111000001111111111111111", 
 "111111111111111000111110000000011111000000111110000111111111111111110000001111111111111111", 
 "111111111111111000111110000000011111000000111110000000000000011111000000001111111111111111", 
 "111111111111111000111110000000011111000000111110000000000000011111000000001111111111111111", 
 "111111111111111000111110000001111111000000111111000000000000011111000000001111111111111111", 
 "111111111111111000111110000001111111000000111111110000000000011111000000001111111111111111", 
 "111111111111111000000000000011111100000000111111110000000000011111000000001111111111111111", 
 "111111111111111000000000001111111000000000111111111111100001111000000000111111111111111111", 
 "111111111111111000000000001111111000000000111111111111100001111000000000111111111111111111", 
 "111111111111111110000000111111100000000000111111111111100001111000000000111111111111111111", 
 "111111111111111110000001111111100000000000111111111110000001111000000000111111111111111111", 
 "111111111111111000000001111100000000000000111111111110000001111000000000111111111111111111", 
 "111111111111111000000111111100000000000011111111111110000011100000000000111111111111111111", 
 "111111111111111000001111111100000000000011111111111110001111100000000111111111111111111111", 
 "111111111111111000001111111100000000000000111111111110001111100000000111111111111111111111", 
 "111111111111111000111111111111111111000000111111111110001111100000000111111111111111111111", 
 "111111111111111000111111111111111111000000111111111110001111100000000111111111111111111111", 
 "111111111111111000000000000000000000000000111111111110000000000000000111111111111111111111", 
 "111111111111111000000000000000000000000000111111111110000000000000111111111111111111111111", 
 "111111111111111000000000000000000000000000111111111110000000000000111111111111111111111111", 
 "111111111111111110000000000000000000000000111111111110000000000000111111111111111111111111", 
 "111111111111111110000000000000000000000000111111111111100000000000111111111111111111111111", 
 "111111111111111111000000000000000000000000111111111111100000000000111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");


Twenty_Eight <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111000000000000000000011111111111111001000000000000100111111111111111111111", 
 "111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111", 
 "111111111111111100000000000000000000000011111111110000000000000000000011111111111111111111", 
 "111111111111111100000011111111111100000011111111000000000000000000000000111111111111111111", 
 "111111111111111100000111111111111100000001111110000001111111111111000000111111111111111111", 
 "111111111111111100011111000000001111100000011110000111110000000011111000000111111111111111", 
 "111111111111111100011111000000001111100000011110000111110000000011111000000111111111111111", 
 "111111111111111100011111000000001111100000011110000111110000000011111000000111111111111111", 
 "111111111111111100011111000000111111100000011110000111110000000011111000000111111111111111", 
 "111111111111111100011111000000111111100000011110000111111100000011111000000111111111111111", 
 "111111111111111100000000000001111110000000011110000111111100000011111000000111111111111111", 
 "111111111111111100000000000111111100000000011110000001111110000111100000000111111111111111", 
 "111111111111111100000000000111111100000000011110000001111111111111000000000111111111111111", 
 "111111111111111100000000000111110000000000011110000001111111111111000000000111111111111111", 
 "111111111111111111000000111111110000000000011110000111110000011111111000000111111111111111", 
 "111111111111111110000000111111100000000000011110000111110000011111111000000111111111111111", 
 "111111111111111100000011111110000000000001111110000111110000000011111000000111111111111111", 
 "111111111111111100000111111110000000000001111110000111110000000011111000000111111111111111", 
 "111111111111111100000111111110000000000001111110000111110000000011111000000111111111111111", 
 "111111111111111100011111111111111111100000011110000001110000000011100000000111111111111111", 
 "111111111111111100011111111111111111100000011110000001111111111111000000000111111111111111", 
 "111111111111111100000000000000000000000000011110000001111111111111000000000111111111111111", 
 "111111111111111100000000000000000000000000011111000000000000000000000000000111111111111111", 
 "111111111111111100000000000000000000000000011111110000000000000000000000000111111111111111", 
 "111111111111111100000000000000000000000000011111110000000000000000000000000111111111111111", 
 "111111111111111111000000000000000000000000011111111110000000000000000000111111111111111111", 
 "111111111111111111000000000000000000000000011111111110000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Twenty_Nine  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111001000000000000100111111111111111111111111111111111111111111111111111111", 
 "111111111111111110000000000000000000011111111111110000000000000000000111111111111111111111", 
 "111111111111111110000000000000000000011111111111110000000000000000000111111111111111111111", 
 "111111111111111000000000000000000000000111111111100000000000000000000011111111111111111111", 
 "111111111111111000001111111111111000000011111110000001000000000000000000111111111111111111", 
 "111111111111111000001111000000111000000001111110000001111111111111000000111111111111111111", 
 "111111111111111000111110000000011111000000111110000001110000000011000000001111111111111111", 
 "111111111111111000111110000000011111000000111110000111100000000011111000001111111111111111", 
 "111111111111111000111110000000011111000000111110000111100000000011111000001111111111111111", 
 "111111111111111000111110000001111111000000111110000111100000000011111000001111111111111111", 
 "111111111111111000111110000001111111000000111110000111100000000011111000001111111111111111", 
 "111111111111111000000000001111111100000000111110000111100000000011111000001111111111111111", 
 "111111111111111000000000001111111000000000111110000001111111111111111000001111111111111111", 
 "111111111111111000000000001111111000000000111110000001111111111111111000001111111111111111", 
 "111111111111111110000001111111100000000000111110000001111111111111111000001111111111111111", 
 "111111111111111110000001111111000000000000111111110000000000000011111000001111111111111111", 
 "111111111111111000000001111100000000000000111111110000000000000011111000001111111111111111", 
 "111111111111111000000111111100000000000011111111111000000000000111000000001111111111111111", 
 "111111111111111000001111111100000000000011111111111110000000011111000000001111111111111111", 
 "111111111111111000001111111110000100000000111111111110000000011111000000001111111111111111", 
 "111111111111111000111111111111111111000000111111111110001111111000000000001111111111111111", 
 "111111111111111000111111111111111111000000111111111110001111111000000000001111111111111111", 
 "111111111111111000000000000000000000000000111111111110001111111000000000001111111111111111", 
 "111111111111111000000000000000000000000000111111111110000000000000000000111111111111111111", 
 "111111111111111000000000000000000000000000111111111110000000000000000000111111111111111111", 
 "111111111111111110000000000000000000000000111111111110000000000000000000111111111111111111", 
 "111111111111111110000000000000000000000000111111111111100000000000000111111111111111111111", 
 "111111111111111111000000000000000000000000111111111111110000000000000111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Thirty       <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111100000000000000000000111111111111100000000000000000011111111111111111111", 
 "111111111111111111100000000000000000000111111111111000000000000000000011111111111111111111", 
 "111111111111111100000000000000000000000001111111110000000000000000000001111111111111111111", 
 "111111111111111100000011111111111110000001111111000000000000000000000000011111111111111111", 
 "111111111111111100000011111111111110000001111111000000111111111111100000011111111111111111", 
 "111111111111111100001111100000000111100000011111000000111000000011100000000111111111111111", 
 "111111111111111100001111100000000111110000001111000011111000000001111100000011111111111111", 
 "111111111111111100000000000000000111110000001111000011111000000001111100000011111111111111", 
 "111111111111111100000000000000000111110000001111000011111000000011111100000011111111111111", 
 "111111111111111100000000000000000111110000001111000011111000001111111100000011111111111111", 
 "111111111111111110000000000000001110000000011111000011111000001111111100000011111111111111", 
 "111111111111111111100000000011111110000000001111000111111000110001111100000111111111111111", 
 "111111111111111111100000000011111110000000001111000011111000110001111100000011111111111111", 
 "111111111111111100000000000000000111000000001111000011111000100001111100000011111111111111", 
 "111111111111111100000000000000000111110000001111000011111110000001111100000011111111111111", 
 "111111111111111100000000000000000111110000001111000011111110000001111100000011111111111111", 
 "111111111111111100001111000000000111110000001111000011111000000001111100000011111111111111", 
 "111111111111111100001111100000000111110000001111000011111000000001111100000011111111111111", 
 "111111111111111100000011100000001111000000011111000011111000000001111100000011111111111111", 
 "111111111111111100000011111111111110000000001111000000111111111111100000000111111111111111", 
 "111111111111111100000011111111111110000000001111000000111111111111100000000011111111111111", 
 "111111111111111110000000000000000000000000001111000000111111111111100000000011111111111111", 
 "111111111111111111100000000000000000000000001111111000000000000000000000000011111111111111", 
 "111111111111111111100000000000000000000000011111111000000000000000000000000011111111111111", 
 "111111111111111111111100000000000000000000111111111000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000001111111111110000000000000000000011111111111111111", 
 "111111111111111111111100000000000000000001111111111111000000000000000000011111111111111111", 
 "111111111111111111111111111111111111111111111111111111000000000000010000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Thirty_One   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111100000000000000000000111111111111111100000000000111111111111111111111111", 
 "111111111111111111100000000000000000000111111111111111100000000000111111111111111111111111", 
 "111111111111111110000000000000000000000001111111111110000000000000001111111111111111111111", 
 "111111111111111100000011111111111110000001111111111100000001111000000111111111111111111111", 
 "111111111111111100000011111111111110000001111111111100000011111000000111111111111111111111", 
 "111111111111111100000011100000000111000000011111111100000011111000000111111111111111111111", 
 "111111111111111100001111100000000111110000001111111100011111111000000111111111111111111111", 
 "111111111111111100000010000000000111110000001111111100000011111000000111111111111111111111", 
 "111111111111111100000000000000000111110000001111111100000011111000000111111111111111111111", 
 "111111111111111100000000000000000111110000001111111100000011111000000111111111111111111111", 
 "111111111111111110000000000000000111000000011111111110000011111000000111111111111111111111", 
 "111111111111111111100000000011111110000000001111111111100011111000000111111111111111111111", 
 "111111111111111111100000000011111110000000001111111111100011111000000111111111111111111111", 
 "111111111111111110000000000000000110000000001111111111100011111000000111111111111111111111", 
 "111111111111111100000000000000000111110000001111111111100011111000000111111111111111111111", 
 "111111111111111100000000000000000111110000001111111111100011111000000111111111111111111111", 
 "111111111111111100001111000000000111110000001111110000000011111000000000111111111111111111", 
 "111111111111111100001111100000000111110000001111110000000011111000000000111111111111111111", 
 "111111111111111100001111100000000111100000001111110000000011111000000000111111111111111111", 
 "111111111111111100000011111111111110000000011111110001111111111111111000000111111111111111", 
 "111111111111111100000011111111111110000000001111110001111111111111110000000111111111111111", 
 "111111111111111100000000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000011111111000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000001111111111100000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000001111111111100000000000000000000000111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Thirty_Two   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111100000000000000000001111111111110000000000000000000111111111111111111111", 
 "111111111111111111100000000000000000000111111111110000000000000000000011111111111111111111", 
 "111111111111111110000000000000000000000001111111000000000000000000000000111111111111111111", 
 "111111111111111100000011111111111110000001111111000000111111111111000000111111111111111111", 
 "111111111111111100000011111111111110000001111111000001111111111111000000011111111111111111", 
 "111111111111111100000011100000000111000000011111000001110000000011100000000111111111111111", 
 "111111111111111100001111100000000111110000001111000111110000000011111000000111111111111111", 
 "111111111111111100001111000000000111110000001111000111110000000011111000000111111111111111", 
 "111111111111111100000000000000000111110000001111000111110000001111111000000111111111111111", 
 "111111111111111100000000000000000111110000001111000111110000001111111000000111111111111111", 
 "111111111111111100000000000000000111100000001111000011110000011111111000000111111111111111", 
 "111111111111111111100000000011111110000000011111000000000001111111000000000111111111111111", 
 "111111111111111111100000000011111110000000001111000000000001111111000000000111111111111111", 
 "111111111111111110000000000000000110000000001111000000000001111100000000000111111111111111", 
 "111111111111111100000000000000000111110000001111110000001111111000000000000111111111111111", 
 "111111111111111100000000000000000111110000001111110000001111111000000000000111111111111111", 
 "111111111111111100001111000000000111110000001111000000111111100000000000011111111111111111", 
 "111111111111111100001111100000000111110000001111000001111111100000000000011111111111111111", 
 "111111111111111100001111100000000111110000001111000001111111100000000000011111111111111111", 
 "111111111111111100000011111111111110000000011111000111111111111111111000000111111111111111", 
 "111111111111111100000011111111111110000000001111000111111111111111111000000111111111111111", 
 "111111111111111100000010000000000000000000001111000001000000000000100000000111111111111111", 
 "111111111111111111100000000000000000000000001111000000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000001111000000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000011111000000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000001111111110000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000001111111110000000000000000000000000111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Thirty_Three <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111100000000000000000000111111111111000000000000000000111111111111111111111", 
 "111111111111111111100000000000000000000111111111110000000000000000000011111111111111111111", 
 "111111111111111100000000000000000000000001111111110000000000000000000011111111111111111111", 
 "111111111111111100000011111111111110000001111111000000000000000000000000111111111111111111", 
 "111111111111111100000011111111111110000000111111000001111111111111000000011111111111111111", 
 "111111111111111100001111100000000111110000011111000001110000000011000000001111111111111111", 
 "111111111111111100001111100000000111110000001111000111110000000011111000000111111111111111", 
 "111111111111111100000000000000000111110000001111000111110000000011111000000111111111111111", 
 "111111111111111100000000000000000111110000001111000000000000000011111000000111111111111111", 
 "111111111111111100000000000000000111110000001111000000000000000011111000000111111111111111", 
 "111111111111111111100000000011111110000000011111000000000000000011111000000111111111111111", 
 "111111111111111111100000000011111110000000001111110000000001111111000000000111111111111111", 
 "111111111111111111100000000011111110000000001111110000000001111111000000000111111111111111", 
 "111111111111111100000000000000000111110000001111110000000001111111000000000111111111111111", 
 "111111111111111100000000000000000111110000001111000000000000000011111000000111111111111111", 
 "111111111111111100000000000000000111110000001111000000000000000011111000000111111111111111", 
 "111111111111111100001111000000000111110000001111000000000000000011111000000111111111111111", 
 "111111111111111100001111100000000111110000001111000111110000000011111000000111111111111111", 
 "111111111111111100000011100000001111000000011111000111110000000011111000000111111111111111", 
 "111111111111111100000011111111111110000000001111000001111111111111000000000111111111111111", 
 "111111111111111100000011111111111110000000001111000001111111111111000000000111111111111111", 
 "111111111111111111000000000000000000000000001111000001111111111111000000000111111111111111", 
 "111111111111111111100000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000011111110000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000001111111111000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000001111111111110000000000000000000011111111111111111", 
 "111111111111111111111100000000000000000001111111111110000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111000000000000100000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Thirty_Four  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111110000000000111111111111111111111", 
 "111111111111111111100000000000000000001111111111111111111100000000000011111111111111111111", 
 "111111111111111111100000000000000000000111111111111111111100000000000011111111111111111111", 
 "111111111111111110000000000000000000000011111111111111110000000000000000111111111111111111", 
 "111111111111111100000011111111111110000001111111111111110000001111000000011111111111111111", 
 "111111111111111100000011111111111110000001111111111111110000011111000000011111111111111111", 
 "111111111111111100000011100000000110000000011111111110000001111111000000011111111111111111", 
 "111111111111111100001111100000000111110000001111111110000001111111000000011111111111111111", 
 "111111111111111100001111000000000111110000001111110000000011111111000000011111111111111111", 
 "111111111111111100000000000000000111110000001111110000001111111111000000011111111111111111", 
 "111111111111111100000000000000000111110000001111110000001111111111000000111111111111111111", 
 "111111111111111100000000000000000111000000011111000000111100011111000000111111111111111111", 
 "111111111111111111100000000011111110000000001111000001111100001111000000111111111111111111", 
 "111111111111111111100000000011111110000000001111000001111100001111000000011111111111111111", 
 "111111111111111110000000000000001110000000001111000111110000001111000000011111111111111111", 
 "111111111111111100000000000000000111110000001111000111110000001111000000011111111111111111", 
 "111111111111111100000000000000000111110000001111000111110000011111100000000111111111111111", 
 "111111111111111100000010000000000111110000001111000111111111111111111000000111111111111111", 
 "111111111111111100001111100000000111110000001111000111111111111111111000000111111111111111", 
 "111111111111111100001111100000000111110000001111000000000000011111000000000111111111111111", 
 "111111111111111100000011111111111110000000011111000000000000001111000000000111111111111111", 
 "111111111111111100000011111111111110000000001111000000000000001111000000000111111111111111", 
 "111111111111111100000010000000000000000000001111100000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000011111111111111111100000000000011111111111111111", 
 "111111111111111111111100000000000000000001111111111111111111100000000000011111111111111111", 
 "111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Thirty_Five  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111100000000000000000000111111111000000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000111111111000000000000000000000000000111111111111111", 
 "111111111111111110000000000000000000000001111111000000000000000000000000000111111111111111", 
 "111111111111111100000011111111111110000001111111000111111111111111111000000111111111111111", 
 "111111111111111100000011111111111110000001111111000111111111111111111000000111111111111111", 
 "111111111111111100000011100000000111000000011111000111110000000000000000000111111111111111", 
 "111111111111111100001111100000000111110000001111000111110000000000000000000111111111111111", 
 "111111111111111100000010000000000111110000001111000111110000000000000000000111111111111111", 
 "111111111111111100000000000000000111110000001111000111111111111111000000000111111111111111", 
 "111111111111111100000000000000000111110000001111000111111111111111000000000111111111111111", 
 "111111111111111110000000000000000111000000011111000000000000000111100000000111111111111111", 
 "111111111111111111100000000011111110000000001111000000000000000011111000000111111111111111", 
 "111111111111111111100000000011111110000000001111000000000000000011111000000111111111111111", 
 "111111111111111110000000000000000110000000001111000000000000000011111000000111111111111111", 
 "111111111111111100000000000000000111110000001111000000000000000011111000000111111111111111", 
 "111111111111111100000000000000000111110000001111000000000000000011111000000111111111111111", 
 "111111111111111100001111000000000111110000001111000111110000000011111000000111111111111111", 
 "111111111111111100001111100000000111110000001111000111110000000011111000000111111111111111", 
 "111111111111111100000111100000000111100000011111000011110000000011110000000111111111111111", 
 "111111111111111100000011111111111110000000001111000001111111111111000000000111111111111111", 
 "111111111111111100000011111111111110000000001111000001111111111111000000000111111111111111", 
 "111111111111111100000000000000000000000000001111000000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000011111111000000000000000000000001111111111111111", 
 "111111111111111111111100000000000000000001111111111110000000000000000000011111111111111111", 
 "111111111111111111111100000000000000000001111111111110000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Thirty_Six   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111110000000000000000000111111111111111000000000000011111111111111111111111", 
 "111111111111111111110000000000000000000011111111111110000000000000011111111111111111111111", 
 "111111111111111111100000000000000000000011111111111110000000000000011111111111111111111111", 
 "111111111111111110000001000000000000000000111111110000000000000000000011111111111111111111", 
 "111111111111111110000001111111111111000000111111110000001111111100000011111111111111111111", 
 "111111111111111110000001110000000011000000001111000000001110000000000011111111111111111111", 
 "111111111111111110000111110000000011111000000111000000111110000000000011111111111111111111", 
 "111111111111111110000111110000000011111000000111000000111110000000000011111111111111111111", 
 "111111111111111110000000000000000011111000000111000001110000000000000011111111111111111111", 
 "111111111111111110000000000000000011111000000111000111110000000000000011111111111111111111", 
 "111111111111111110000000000000000011111000000111000111110000000000000011111111111111111111", 
 "111111111111111111110000000001111111000000001111000111111111111111100000011111111111111111", 
 "111111111111111111110000000001111111000000000111000111111111111111000000011111111111111111", 
 "111111111111111111000000000000000111000000000111000111111000000111100000001111111111111111", 
 "111111111111111110000000000000000011111000000111000111110000000011111000000111111111111111", 
 "111111111111111110000000000000000011111000000111000111110000000001111000000111111111111111", 
 "111111111111111110000000000000000011111000000111000111110000000001111000000111111111111111", 
 "111111111111111110000111110000000011111000000111000111110000000001111000000111111111111111", 
 "111111111111111110000111110000000011111000000111000111110000000001111000000111111111111111", 
 "111111111111111110000001111111111111000000001111000001111111111111100000000111111111111111", 
 "111111111111111110000001111111111111000000000111000000111111111111000000000111111111111111", 
 "111111111111111110000001111111111111000000000111000000111111111111000000000111111111111111", 
 "111111111111111111110000000000000000000000000111110000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000000111110000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000001111111000000000000000000000000111111111111111", 
 "111111111111111111111110000000000000000000111111111110000000000000000000011111111111111111", 
 "111111111111111111111110000000000000000000111111111110000000000000000000111111111111111111", 
 "111111111111111111111111000000000000100001111111111111000111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Thirty_Seven <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111000000000000000000000000111111111111111111", 
 "111111111111111111100000000000000000001111111111000000000000000000000000111111111111111111", 
 "111111111111111111100000000000000000000111111111000000000000000000000000011111111111111111", 
 "111111111111111110000000000000000000000011111111000000000000000000100000000111111111111111", 
 "111111111111111100000011111111111110000001111111000111111111111111111000000111111111111111", 
 "111111111111111100000011111111111110000001111111000111111111111111111000000111111111111111", 
 "111111111111111100000011100000000110000000011111000000000000001111000000000111111111111111", 
 "111111111111111100001111100000000111110000001111000000000000001111000000000111111111111111", 
 "111111111111111100001111000000000111110000001111000000000000001111000000000111111111111111", 
 "111111111111111100000000000000000111110000001111110000000000001111000000000111111111111111", 
 "111111111111111100000000000000000111110000001111110000000000011111000000000111111111111111", 
 "111111111111111100000000000000000111000000011111111111110001111100000000011111111111111111", 
 "111111111111111111100000000011111110000000001111111111110001111000000000111111111111111111", 
 "111111111111111111100000000011111110000000001111111111110001111000000000011111111111111111", 
 "111111111111111110000000000000001110000000001111111110000001111000000000011111111111111111", 
 "111111111111111100000000000000000111110000001111111110000001111000000000111111111111111111", 
 "111111111111111100000000000000000111110000001111111110000001100000000000111111111111111111", 
 "111111111111111100000010000000000111110000001111111110001111100000000011111111111111111111", 
 "111111111111111100001111100000000111110000001111111110001111100000000011111111111111111111", 
 "111111111111111100001111100000000111110000001111111110001111100000000011111111111111111111", 
 "111111111111111100000011111111111110000000011111111110001111100000000011111111111111111111", 
 "111111111111111100000011111111111110000000001111111110000000000000000111111111111111111111", 
 "111111111111111100000010000000000000000000001111111110000000000000011111111111111111111111", 
 "111111111111111111100000000000000000000000001111111110000000000000011111111111111111111111", 
 "111111111111111111100000000000000000000000001111111110000000000000011111111111111111111111", 
 "111111111111111111110000000000000000000000011111111111110000000000011111111111111111111111", 
 "111111111111111111111100000000000000000001111111111111110000000000011111111111111111111111", 
 "111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Thirty_Eight <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111001000000000000100111111111111001000000000000100111111111111111111111", 
 "111111111111111111110000000000000000000011111111110000000000000000000011111111111111111111", 
 "111111111111111111110000000000000000000011111111110000000000000000000011111111111111111111", 
 "111111111111111110000000000000000000000000111111000000000000000000000000111111111111111111", 
 "111111111111111110000001111111111111000000111111000000111111111111000000011111111111111111", 
 "111111111111111110000001111111111111000000111111000011110000000011111000000111111111111111", 
 "111111111111111110000111110000000011111000000111000111110000000001111000000111111111111111", 
 "111111111111111110000111110000000011111000000111000111110000000001111000000111111111111111", 
 "111111111111111110000000000000000011111000000111000111110000000001111000000111111111111111", 
 "111111111111111110000000000000000011111000000111000111111100000001111000000111111111111111", 
 "111111111111111110000000000000000011111000000111000111111110000011111000000111111111111111", 
 "111111111111111111000000000000000111000000001111000001111110000011100000000111111111111111", 
 "111111111111111111110000000001111111000000000111000000111111111111000000000111111111111111", 
 "111111111111111111110000000001111111000000000111000000111111111111000000000111111111111111", 
 "111111111111111110000000000000000011110000000111000011110000001111111000000111111111111111", 
 "111111111111111110000000000000000011111000000111000111110000001111111000000111111111111111", 
 "111111111111111110000000000000000011111000000111000111110000000011111000000111111111111111", 
 "111111111111111110000111110000000011111000000111000111110000000001111000000111111111111111", 
 "111111111111111110000111110000000011111000000111000111110000000001111000000111111111111111", 
 "111111111111111110000001110000000011100000001111000001110000000011100000000111111111111111", 
 "111111111111111110000001111111111111000000000111000000111111111111000000000111111111111111", 
 "111111111111111110000001111111111111000000000111000000111111111111000000000111111111111111", 
 "111111111111111111000000000000000000000000000111000000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000000111110000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000001111111000000000000000000000000111111111111111", 
 "111111111111111111111110000000000000000000111111111110000000000000000000011111111111111111", 
 "111111111111111111111110000000000000000000111111111110000000000000000000011111111111111111", 
 "111111111111111111111110000000000000000000111111111111000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



Thirty_Nine  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111100000000000000000001111111111110000000000000000000111111111111111111111", 
 "111111111111111111100000000000000000000111111111110000000000000000000011111111111111111111", 
 "111111111111111111000000000000000000000111111111100000000000000000000011111111111111111111", 
 "111111111111111100000010000000000000000001111111000000000000000000000000111111111111111111", 
 "111111111111111100000011111111111110000001111111000001111111111111000000011111111111111111", 
 "111111111111111100000011100000000110000000011111000001110000000011100000001111111111111111", 
 "111111111111111100001111100000000111110000001111000111110000000011111000000111111111111111", 
 "111111111111111100001111000000000111110000001111000111110000000011111000000111111111111111", 
 "111111111111111100000000000000000111110000001111000111110000000011111000000111111111111111", 
 "111111111111111100000000000000000111110000001111000111110000000011111000000111111111111111", 
 "111111111111111100000000000000000111110000001111000111110000000011111000000111111111111111", 
 "111111111111111111100000000011111110000000011111000001111111111111111000000111111111111111", 
 "111111111111111111100000000011111110000000001111000001111111111111111000000111111111111111", 
 "111111111111111111000000000011111110000000001111000000111111111111111000000111111111111111", 
 "111111111111111100000000000000000111110000001111110000000000000011111000000111111111111111", 
 "111111111111111100000000000000000111110000001111110000000000000011111000000111111111111111", 
 "111111111111111100000000000000000111110000001111111000000000000011000000000111111111111111", 
 "111111111111111100001111100000000111110000001111111110000000001111000000000111111111111111", 
 "111111111111111100001111100000000111110000001111111110000000011111000000000111111111111111", 
 "111111111111111100000011111111111110000000011111111110001111111100000000000111111111111111", 
 "111111111111111100000011111111111110000000001111111110001111111100000000000111111111111111", 
 "111111111111111100000011111111111110000000001111111110001111111000000000000111111111111111", 
 "111111111111111111100000000000000000000000001111111110000000000000000000011111111111111111", 
 "111111111111111111100000000000000000000000001111111110000000000000000000111111111111111111", 
 "111111111111111111100000000000000000000000011111111110000000000000000000111111111111111111", 
 "111111111111111111111100000000000000000001111111111111110000000000000011111111111111111111", 
 "111111111111111111111100000000000000000001111111111111110000000000000111111111111111111111", 
 "111111111111111111111110000000000011100011111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



forty        <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111100000000001111111111111000000000000000000111111111111111111111", 
 "111111111111111111111111111000000000000111111111110000000000000000000011111111111111111111", 
 "111111111111111111111111111000000000000111111111110000000000000000000011111111111111111111", 
 "111111111111111111111111100000000000000001111111000000000000000000000000111111111111111111", 
 "111111111111111111111111100000111110000001111111000001111111111111000000011111111111111111", 
 "111111111111111111111110000000111110000001111111000001110000000111000000001111111111111111", 
 "111111111111111111111100000011111110000001111111000111110000000011111000000111111111111111", 
 "111111111111111111111100000011111110000001111111000111110000000011111000000111111111111111", 
 "111111111111111111100000000111111110000001111111000111110000000011111000000111111111111111", 
 "111111111111111111100000011111111110000001111111000111110000001111111000000111111111111111", 
 "111111111111111111100000011111111110000001111111000111110000001111111000000111111111111111", 
 "111111111111111110000011111000111110000001111111000111110001100011111000000111111111111111", 
 "111111111111111100000011111000111110000001111111000111110001100011111000000111111111111111", 
 "111111111111111100000011110000111110000001111111000111110001000011111000000111111111111111", 
 "111111111111111100001111100000111110000001111111000111111100000011111000000111111111111111", 
 "111111111111111100001111100000111110000001111111000111111100000011111000000111111111111111", 
 "111111111111111100001111100000111111000000011111000111110000000011111000000111111111111111", 
 "111111111111111100001111111111111111110000001111000111110000000011111000000111111111111111", 
 "111111111111111100001111111111111111110000001111000111110000000011111000000111111111111111", 
 "111111111111111110000000000000111110000000001111000001111111111111100000000111111111111111", 
 "111111111111111100000000000000111110000000001111000001111111111111000000000111111111111111", 
 "111111111111111100000000000000011110000000001111000000111111111111000000000111111111111111", 
 "111111111111111111100000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000011111110000000000000000000000000111111111111111", 
 "111111111111111111111111111111000000000000111111111110000000000000000000011111111111111111", 
 "111111111111111111111111111111000000000001111111111110000000000000000000011111111111111111", 
 "111111111111111111111111111111000000000001111111111111000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");


forty_one    <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111000000000000111111111111111111111111", 
 "111111111111111111111111111000000000000111111111111111000000000000111111111111111111111111", 
 "111111111111111111111111111000000000000111111111111100000000000000001111111111111111111111", 
 "111111111111111111111111100000000000000001111111111100000011110000001111111111111111111111", 
 "111111111111111111111111100000111110000001111111111100000011110000001111111111111111111111", 
 "111111111111111111111111000000111110000001111111111100000111110000001111111111111111111111", 
 "111111111111111111111100000001111110000001111111111100011111110000001111111111111111111111", 
 "111111111111111111111100000011111110000001111111111100000111110000001111111111111111111111", 
 "111111111111111111110000000011111110000001111111111100000011110000001111111111111111111111", 
 "111111111111111111100000011111111110000001111111111100000011110000001111111111111111111111", 
 "111111111111111111100000011111111110000001111111111100000011110000001111111111111111111111", 
 "111111111111111110000011111100111110000001111111111111000011110000001111111111111111111111", 
 "111111111111111100000011111000111110000001111111111111000011110000001111111111111111111111", 
 "111111111111111100000011111000111110000001111111111111000011110000001111111111111111111111", 
 "111111111111111100000111100000111110000001111111111111000011110000001111111111111111111111", 
 "111111111111111100001111100000111110000001111111111111000011110000001111111111111111111111", 
 "111111111111111100001111100000111110000000011111100000000011110000000001111111111111111111", 
 "111111111111111100001111111111111111110000001111100000000011110000000001111111111111111111", 
 "111111111111111100001111111111111111110000001111100000000011111000000001111111111111111111", 
 "111111111111111100000000000000111111000000001111100011111111111111110000001111111111111111", 
 "111111111111111100000000000000111110000000001111100001111111111111110000001111111111111111", 
 "111111111111111100000000000000111110000000001111100000000000000000000000001111111111111111", 
 "111111111111111110000000000000000000000000001111100000000000000000000000001111111111111111", 
 "111111111111111111100000000000000000000000001111100000000000000000000000001111111111111111", 
 "111111111111111111100000000000000000000000001111110000000000000000000000001111111111111111", 
 "111111111111111111111111111111000000000000111111111100000000000000000000001111111111111111", 
 "111111111111111111111111111111000000000001111111111100000000000000000000001111111111111111", 
 "111111111111111111111111111111000000000001111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");


forty_two    <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111100000000000011111111111000000000000000000011111111111111111111", 
 "111111111111111111111111111100000000000011111111110000000000000000000011111111111111111111", 
 "111111111111111111111111110000000000000000111111000000000000000000000000111111111111111111", 
 "111111111111111111111111110000001111000000111111000000111111111111000000011111111111111111", 
 "111111111111111111111111110000011111000000111111000000111111111111100000011111111111111111", 
 "111111111111111111111110000000011111000000111111000001110000000011100000000111111111111111", 
 "111111111111111111111110000001111111000000111111000111110000000001111000000111111111111111", 
 "111111111111111111111110000001111111000000111111000111110000000001111000000111111111111111", 
 "111111111111111111110000001111111111000000111111000111110000001111111000000111111111111111", 
 "111111111111111111110000001111111111000000111111000111110000001111111000000111111111111111", 
 "111111111111111111100000001111111111000000111111000011110000001111111000000111111111111111", 
 "111111111111111110000001111100011111000000111111000000000001111111100000000111111111111111", 
 "111111111111111110000001111100011111000000111111000000000001111111100000000111111111111111", 
 "111111111111111110000001110000011111000000111111000000000001111100000000000111111111111111", 
 "111111111111111110000111110000011111000000111111110000000111111100000000000111111111111111", 
 "111111111111111110000111110000011111000000011111110000001111111000000000000111111111111111", 
 "111111111111111110000111111111111111110000000111000000111111100000000000011111111111111111", 
 "111111111111111110000111111111111111111000000111000000111111100000000000011111111111111111", 
 "111111111111111110000111111111111111111000000111000000111111100000000000011111111111111111", 
 "111111111111111110000000000000011111000000000111000111111111111111111000000111111111111111", 
 "111111111111111110000000000000011111000000000111000111111111111111111000000111111111111111", 
 "111111111111111111000000000000000000000000000111000001000000000000110000000111111111111111", 
 "111111111111111111110000000000000000000000000111000000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000000111000000000000000000000000000111111111111111", 
 "111111111111111111111001000000000000000000001111000000000000000000000000000111111111111111", 
 "111111111111111111111111111111100000000000111111110000000000000000000000000111111111111111", 
 "111111111111111111111111111111100000000000111111111000000000000000000000000111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");


forty_three  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111110000000000111111111111000000000000000000011111111111111111111", 
 "111111111111111111111111111100000000000011111111110000000000000000000011111111111111111111", 
 "111111111111111111111111111100000000000011111111110000000000000000000011111111111111111111", 
 "111111111111111111111111110000000000000000111111000000000000000000000000011111111111111111", 
 "111111111111111111111111110000011111000000111111000000111111111111100000011111111111111111", 
 "111111111111111111111110000000011111000000111111000000110000000011100000000111111111111111", 
 "111111111111111111111110000001111111000000111111000111110000000001111000000111111111111111", 
 "111111111111111111111110000001111111000000111111000011110000000001111000000111111111111111", 
 "111111111111111111110000000011111111000000111111000000000000000001111000000111111111111111", 
 "111111111111111111110000001111111111000000111111000000000000000001111000000111111111111111", 
 "111111111111111111110000001111111111000000111111000000000000000001111000000111111111111111", 
 "111111111111111110000001111100011111000000111111111000000001111111100000000111111111111111", 
 "111111111111111110000001111100011111000000111111110000000001111111100000000111111111111111", 
 "111111111111111110000001111100011111000000111111110000000000111111100000000111111111111111", 
 "111111111111111110000111110000011111000000111111000000000000000001111000000111111111111111", 
 "111111111111111110000111110000011111000000011111000000000000000001111000000111111111111111", 
 "111111111111111110000111110000011111100000001111000000000000000001111000000111111111111111", 
 "111111111111111110000111111111111111111000000111000111110000000001111000000111111111111111", 
 "111111111111111110000111111111111111111000000111000111110000000001111000000111111111111111", 
 "111111111111111110000000000000011111000000000111000000111111111111100000000111111111111111", 
 "111111111111111110000000000000011111000000000111000000111111111111100000000111111111111111", 
 "111111111111111110000000000000011111000000000111000000111111111111100000000111111111111111", 
 "111111111111111111110000000000000000000000000111110000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000000111110000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000001111111000000000000000000000000111111111111111", 
 "111111111111111111111111111111100000000000111111111110000000000000000000011111111111111111", 
 "111111111111111111111111111111100000000000111111111110000000000000000000011111111111111111", 
 "111111111111111111111111111111100000000000111111111111000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");


forty_four   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111110000000000111111111111111111110000000000011111111111111111111", 
 "111111111111111111111111111100000000000011111111111111111110000000000011111111111111111111", 
 "111111111111111111111111111100000000000011111111111111111100000000000011111111111111111111", 
 "111111111111111111111111110000000000000000111111111111110000000000000000011111111111111111", 
 "111111111111111111111111110000011111000000111111111111110000001111100000011111111111111111", 
 "111111111111111111111111100000011111000000111111111111110000001111100000011111111111111111", 
 "111111111111111111111110000001111111000000111111111110000001111111100000011111111111111111", 
 "111111111111111111111110000001111111000000111111111110000001111111100000011111111111111111", 
 "111111111111111111110000000011111111000000111111111000000001111111100000011111111111111111", 
 "111111111111111111110000001111111111000000111111110000000111111111100000011111111111111111", 
 "111111111111111111110000001111111111000000111111110000001111111111100000011111111111111111", 
 "111111111111111111000001111100011111000000111111000000111110001111100000011111111111111111", 
 "111111111111111110000001111100011111000000111111000000111110001111100000011111111111111111", 
 "111111111111111110000001111100011111000000111111000000111100001111100000011111111111111111", 
 "111111111111111110000111110000011111000000111111000111110000001111100000011111111111111111", 
 "111111111111111110000111110000011111000000111111000111110000001111100000011111111111111111", 
 "111111111111111110000111110000011111100000001111000111110000011111100000000111111111111111", 
 "111111111111111110000111111111111111111000000111000111111111111111111000000111111111111111", 
 "111111111111111110000111111111111111111000000111000111111111111111111000000111111111111111", 
 "111111111111111110000000000000011111000000000111000000000000001111100000000111111111111111", 
 "111111111111111110000000000000011111000000000111000000000000001111100000000111111111111111", 
 "111111111111111110000000000000001111000000000111000000000000001111000000000111111111111111", 
 "111111111111111111100000000000000000000000000111110000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000000111110000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000001111111000000000000000000000000111111111111111", 
 "111111111111111111111111111111100000000000111111111111111111100000000000011111111111111111", 
 "111111111111111111111111111111100000000000111111111111111111100000000000011111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");


forty_five   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111000000000000111111110000000000000000000000000001111111111111111", 
 "111111111111111111111111111000000000000111111110000000000000000000000000001111111111111111", 
 "111111111111111111111111100000000000000001111110000000000000000000000000001111111111111111", 
 "111111111111111111111111100000011110000001111110000111111111111111110000001111111111111111", 
 "111111111111111111111111100000111110000001111110001111111111111111110000001111111111111111", 
 "111111111111111111111100000000111110000001111110001111100000000000000000001111111111111111", 
 "111111111111111111111100000011111110000001111110001111100000000000000000001111111111111111", 
 "111111111111111111110000000011111110000001111110001111100000000000000000001111111111111111", 
 "111111111111111111100000011111111110000001111110001111111111111110000000001111111111111111", 
 "111111111111111111100000011111111110000001111110001111111111111111000000001111111111111111", 
 "111111111111111110000000011100111110000001111110000000000000000111000000001111111111111111", 
 "111111111111111100000011111000111110000001111110000000000000000011110000001111111111111111", 
 "111111111111111100000011111000111110000001111110000000000000000011110000001111111111111111", 
 "111111111111111100000011100000111110000001111110000000000000000011110000001111111111111111", 
 "111111111111111100001111100000111110000001111110000000000000000011110000001111111111111111", 
 "111111111111111100001111100000111110000000111110000000000000000011110000001111111111111111", 
 "111111111111111100001111111111111111100000001110000111100000000011110000001111111111111111", 
 "111111111111111100001111111111111111110000001110001111100000000011110000001111111111111111", 
 "111111111111111100000111111111111111100000001110000111100000000111110000001111111111111111", 
 "111111111111111100000000000000111110000000001110000001111111111111000000001111111111111111", 
 "111111111111111100000000000000111110000000001110000001111111111111000000001111111111111111", 
 "111111111111111110000000000000000000000000001110000000000000000000000000001111111111111111", 
 "111111111111111111100000000000000000000000001111100000000000000000000000001111111111111111", 
 "111111111111111111100000000000000000000000001111100000000000000000000000001111111111111111", 
 "111111111111111111110010000000000000000000011111111000000000000000000000011111111111111111", 
 "111111111111111111111111111111000000000001111111111100000000000000000000111111111111111111", 
 "111111111111111111111111111111000000000001111111111100000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");


forty_six    <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111100000000001111111111111100000000000001111111111111111111111111", 
 "111111111111111111111111111000000000000111111111111000000000000001111111111111111111111111", 
 "111111111111111111111111110000000000000111111111111000000000000000111111111111111111111111", 
 "111111111111111111111111100000000000000001111111100000000000000000001111111111111111111111", 
 "111111111111111111111111100000111110000001111111100000011111110000001111111111111111111111", 
 "111111111111111111111100000000111110000001111110000000011000000000001111111111111111111111", 
 "111111111111111111111100000011111110000001111100000011111000000000001111111111111111111111", 
 "111111111111111111111100000011111110000001111100000011111000000000001111111111111111111111", 
 "111111111111111111100000000111111110000001111100000111000000000000001111111111111111111111", 
 "111111111111111111100000011111111110000001111100001111000000000000001111111111111111111111", 
 "111111111111111111100000011111111110000001111100001111000000000000001111111111111111111111", 
 "111111111111111100000011111000111110000001111100011111111111111110000001111111111111111111", 
 "111111111111111100000011111000111110000001111100001111111111111110000001111111111111111111", 
 "111111111111111100000011100000111110000001111100001111100000001110000000011111111111111111", 
 "111111111111111100001111100000111110000001111100001111000000000111110000011111111111111111", 
 "111111111111111100001111100000111110000001111100001111000000000111110000011111111111111111", 
 "111111111111111100001111100000111111000000011100001111000000000111110000011111111111111111", 
 "111111111111111100001111111111111111110000001100001111000000000111110000011111111111111111", 
 "111111111111111100001111111111111111110000001100001111000000000111110000011111111111111111", 
 "111111111111111110000000000000111110000000001100000011111111111110000000011111111111111111", 
 "111111111111111100000000000000111110000000001100000011111111111110000000011111111111111111", 
 "111111111111111100000000000000011110000000001100000011111111111110000000011111111111111111", 
 "111111111111111111100000000000000000000000001111100000000000000000000000011111111111111111", 
 "111111111111111111100000000000000000000000001111100000000000000000000000011111111111111111", 
 "111111111111111111100000000000000000000000011111100000000000000000000000011111111111111111", 
 "111111111111111111111111111111000000000001111111111000000000000000000001111111111111111111", 
 "111111111111111111111111111111000000000001111111111000000000000000000001111111111111111111", 
 "111111111111111111111111111111100001000011111111111110001111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");


forty_seven  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111100000000001111111110000000000000000000000001111111111111111111", 
 "111111111111111111111111111000000000000111111110000000000000000000000000111111111111111111", 
 "111111111111111111111111111000000000000111111110000000000000000000000000111111111111111111", 
 "111111111111111111111111100000000000000001111110000000000000000000000000001111111111111111", 
 "111111111111111111111111100000111110000001111110001111111111111111110000001111111111111111", 
 "111111111111111111111111000000111110000001111110000111111111111111110000001111111111111111", 
 "111111111111111111111100000011111110000001111110000000000000011111000000001111111111111111", 
 "111111111111111111111100000011111110000001111110000000000000011111000000001111111111111111", 
 "111111111111111111100000000111111110000001111110000000000000011111000000001111111111111111", 
 "111111111111111111100000011111111110000001111111100000000000011111000000001111111111111111", 
 "111111111111111111100000011111111110000001111111110000000000011110000000001111111111111111", 
 "111111111111111110000011111000111110000001111111111111100001111000000000111111111111111111", 
 "111111111111111100000011111000111110000001111111111111100011111000000000111111111111111111", 
 "111111111111111100000011111000111110000001111111111111100011111000000000111111111111111111", 
 "111111111111111100001111100000111110000001111111111100000011111000000000111111111111111111", 
 "111111111111111100001111100000111110000001111111111100000011111000000000111111111111111111", 
 "111111111111111100001111100000111111000000011111111100000011100000000001111111111111111111", 
 "111111111111111100001111111111111111110000001111111100001111000000000111111111111111111111", 
 "111111111111111100001111111111111111110000001111111100011111000000000111111111111111111111", 
 "111111111111111100000000000000111110000000001111111100011111000000000111111111111111111111", 
 "111111111111111100000000000000111110000000001111111100001111000000000111111111111111111111", 
 "111111111111111100000000000000011110000000001111111100000000000000000111111111111111111111", 
 "111111111111111111000000000000000000000000001111111100000000000000111111111111111111111111", 
 "111111111111111111100000000000000000000000001111111100000000000000111111111111111111111111", 
 "111111111111111111100000000000000000000000011111111110000000000000111111111111111111111111", 
 "111111111111111111111111111111000000000001111111111111100000000000111111111111111111111111", 
 "111111111111111111111111111111000000000001111111111111100000000000111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



forty_eight  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111100000001001111111111110110000000000001001111111111111111111111", 
 "111111111111111111111111111000000000000111111111100000000000000000001111111111111111111111", 
 "111111111111111111111111111000000000000111111111100000000000000000001111111111111111111111", 
 "111111111111111111111111100000000000000001111100000000000000000000000001111111111111111111", 
 "111111111111111111111111100000011110000001111100000011111111111110000001111111111111111111", 
 "111111111111111111111111100000111110000001111100001111000000000111100000011111111111111111", 
 "111111111111111111111100000011111110000001111100001111000000000111110000011111111111111111", 
 "111111111111111111111100000011111110000001111100001111000000000111110000011111111111111111", 
 "111111111111111111100000000011111110000001111100001111100000000111110000011111111111111111", 
 "111111111111111111100000011111111110000001111100001111111000000111110000011111111111111111", 
 "111111111111111111100000011111111110000001111100001111111000000111110000011111111111111111", 
 "111111111111111110000000011100111110000001111100000011111100001110000000011111111111111111", 
 "111111111111111100000011111000111110000001111100000011111111111110000000011111111111111111", 
 "111111111111111100000011111000111110000001111100000011111111111110000000011111111111111111", 
 "111111111111111100000111100000111110000001111100001111000000111111100000011111111111111111", 
 "111111111111111100001111100000111110000001111100001111000000111111110000011111111111111111", 
 "111111111111111100001111100000111110000000011100001111000000001111110000011111111111111111", 
 "111111111111111100001111111111111111110000001100001111000000000111110000011111111111111111", 
 "111111111111111100001111111111111111110000001100001111000000000111110000011111111111111111", 
 "111111111111111100000000000000111111000000001100000111100000001110000000011111111111111111", 
 "111111111111111100000000000000111110000000001100000011111111111110000000011111111111111111", 
 "111111111111111100000000000000111110000000001100000011111111111110000000011111111111111111", 
 "111111111111111110000000000000000000000000001100000000000000000000000000011111111111111111", 
 "111111111111111111100000000000000000000000001111100000000000000000000000011111111111111111", 
 "111111111111111111100000000000000000000000001111100000000000000000000000011111111111111111", 
 "111111111111111111111111111111000000000000111111111000000000000000000001111111111111111111", 
 "111111111111111111111111111111000000000001111111111000000000000000000001111111111111111111", 
 "111111111111111111111111111111000000000001111111111100000000000000000001111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



forty_nine   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111000000000011111111111100000000000000000001111111111111111111111", 
 "111111111111111111111111110000000000001111111111000000000000000000001111111111111111111111", 
 "111111111111111111111111110000000000001111111111000000000000000000001111111111111111111111", 
 "111111111111111111111111000000000000000011111100000000000000000000000001111111111111111111", 
 "111111111111111111111111000001111100000011111100000011111111111110000001111111111111111111", 
 "111111111111111111111000000001111100000011111100000111000000001110000000011111111111111111", 
 "111111111111111111111000000111111100000011111100011111000000000111100000011111111111111111", 
 "111111111111111111111000000111111100000011111100011111000000000111100000011111111111111111", 
 "111111111111111111000000111111111100000011111100011111000000000111100000011111111111111111", 
 "111111111111111111000000111111111100000011111100011111000000000111100000011111111111111111", 
 "111111111111111111000000111111111100000011111100011111000000000111100000011111111111111111", 
 "111111111111111000000111110001111100000011111100000011111111111111100000011111111111111111", 
 "111111111111111000000111110001111100000011111100000011111111111111100000011111111111111111", 
 "111111111111111000000111110001111100000011111100000011111111111111100000011111111111111111", 
 "111111111111111000011111000001111100000011111111000000000000000111100000011111111111111111", 
 "111111111111111000011111000001111100000001111111100000000000000111100000011111111111111111", 
 "111111111111111000011111000001111110000000011111100000000000001110000000011111111111111111", 
 "111111111111111000011111111111111111100000011111111000000000111110000000011111111111111111", 
 "111111111111111000011111111111111111100000011111111000000000111100000000011111111111111111", 
 "111111111111111000000000000001111100000000011111111000011111110000000000011111111111111111", 
 "111111111111111000000000000001111100000000011111111000011111110000000000011111111111111111", 
 "111111111111111000000000000000111100000000011111111000011111110000000000011111111111111111", 
 "111111111111111111000000000000000000000000011111111000000000000000000001111111111111111111", 
 "111111111111111111000000000000000000000000011111111000000000000000000001111111111111111111", 
 "111111111111111111100000000000000000000000111111111100000000000000000011111111111111111111", 
 "111111111111111111111111111110000000000011111111111111000000000000001111111111111111111111", 
 "111111111111111111111111111110000000000011111111111111000000000000001111111111111111111111", 
 "111111111111111111111111111111000111000111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



fifty        <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111000000000000000000000000000111111110000000000000000000111111111111111111111", 
 "111111111111111000000000000000000000000000111111110000000000000000000111111111111111111111", 
 "111111111111111000000000000000000000000000111111100000000000000000000111111111111111111111", 
 "111111111111111000011111111111111111100000111110000000000000000000000000111111111111111111", 
 "111111111111111000011111111111111111000000111110000001111111111111000000111111111111111111", 
 "111111111111111000011110000000000000000000111110000001110000000111000000001111111111111111", 
 "111111111111111000011110000000000000000000111110001111100000000011110000001111111111111111", 
 "111111111111111000011111000000000000000000111110001111100000000011111000001111111111111111", 
 "111111111111111000011111111111111100000000111110001111100000000111111000001111111111111111", 
 "111111111111111000011111111111111100000000111110001111100000011111111000001111111111111111", 
 "111111111111111000000000000000001110000000111110001111100000011111111000001111111111111111", 
 "111111111111111000000000000000001111100000111110001111100011000011111000001111111111111111", 
 "111111111111111000000000000000001111100000111110001111100001000011111000001111111111111111", 
 "111111111111111000000000000000001111100000111110001111100001000011111000001111111111111111", 
 "111111111111111000000000000000001111100000111110001111111100000011111000001111111111111111", 
 "111111111111111000000000000000001111100000111110001111111100000011111000001111111111111111", 
 "111111111111111000011110000000001111100000111110001111110000000011111000001111111111111111", 
 "111111111111111000011110000000001111100000111110001111100000000011111000001111111111111111", 
 "111111111111111000000111000000011100000000111110001111100000000011111000001111111111111111", 
 "111111111111111000000111111111111100000000111110000001111111111111000000001111111111111111", 
 "111111111111111000000111111111111100000000111110000001111111111111000000001111111111111111", 
 "111111111111111000000000000000000000000000111110000001111111111111000000001111111111111111", 
 "111111111111111111000000000000000000000000111111100000000000000000000000001111111111111111", 
 "111111111111111111000000000000000000000000111111110000000000000000000000001111111111111111", 
 "111111111111111111110000000000000000000011111111110000000000000000000000001111111111111111", 
 "111111111111111111111000000000000000000011111111111100000000000000000000111111111111111111", 
 "111111111111111111111000000000000000000011111111111100000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



fifty_one    <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111100000000000111111111111111111111111", 
 "111111111111111100000000000000000000000000011111111111100000000000111111111111111111111111", 
 "111111111111111100000000000000000000000000011111111110000000000000001111111111111111111111", 
 "111111111111111100000000000000000000000000011111111100000011111000000111111111111111111111", 
 "111111111111111100001111111111111111110000011111111100000011111000000111111111111111111111", 
 "111111111111111100001111111111111111100000011111111100000011111000000111111111111111111111", 
 "111111111111111100001111000000000000000000011111111100011111111000000111111111111111111111", 
 "111111111111111100001111000000000000000000011111111100010111111000000111111111111111111111", 
 "111111111111111100001111100000000000000000011111111100000011111000000111111111111111111111", 
 "111111111111111100001111111111111110000000011111111100000011111000000111111111111111111111", 
 "111111111111111100001111111111111110000000011111111110000011111000000111111111111111111111", 
 "111111111111111100000000000000000111100000011111111111100011111000000111111111111111111111", 
 "111111111111111100000000000000000111110000011111111111100011111000000111111111111111111111", 
 "111111111111111100000000000000000111110000011111111111100011111000000111111111111111111111", 
 "111111111111111100000000000000000111110000011111111111100011111000000111111111111111111111", 
 "111111111111111100000000000000000111110000011111111111100011111000000111111111111111111111", 
 "111111111111111100000000000000000111110000011111110000000011111000000000111111111111111111", 
 "111111111111111100001111000000000111110000011111100000000011111000000000111111111111111111", 
 "111111111111111100001111000000000111110000011111100000000011111000000000111111111111111111", 
 "111111111111111100000111100000000111000000011111100001111111111111110000001111111111111111", 
 "111111111111111100000011111111111110000000011111100001111111111111110000001111111111111111", 
 "111111111111111100000011111111111110000000011111100000000000000000000000001111111111111111", 
 "111111111111111110000000000000000000000000011111100000000000000000000000001111111111111111", 
 "111111111111111111100000000000000000000000011111100000000000000000000000001111111111111111", 
 "111111111111111111100000000000000000000000011111110000000000000000000000001111111111111111", 
 "111111111111111111111000000000000000000001111111111100000000000000000000001111111111111111", 
 "111111111111111111111100000000000000000001111111111100000000000000000000001111111111111111", 
 "111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




fifty_two    <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111100000000000000000000000000011111110000000000000000000111111111111111111111", 
 "111111111111111100000000000000000000000000011111110000000000000000000111111111111111111111", 
 "111111111111111100000000000000000000000000011111000000000000000000000000111111111111111111", 
 "111111111111111100001111111111111111100000011110000001111111111111000000111111111111111111", 
 "111111111111111100001111111111111111110000011110000001111111111111000000111111111111111111", 
 "111111111111111100001111000000000000000000011110000001110000000011100000001111111111111111", 
 "111111111111111100001111000000000000000000011110000111110000000011111000000111111111111111", 
 "111111111111111100001111000000000000000000011110000111110000000011111000000111111111111111", 
 "111111111111111100001111111111111100000000011110000111110000001111111000000111111111111111", 
 "111111111111111100001111111111111110000000011110000111110000011111111000000111111111111111", 
 "111111111111111100001111111111111110000000011110000111100000011111110000001111111111111111", 
 "111111111111111100000000000000000111110000011110000000000001111111000000001111111111111111", 
 "111111111111111100000000000000000111110000011110000000000001111111000000000111111111111111", 
 "111111111111111100000000000000000111110000011111000000000011111100000000000111111111111111", 
 "111111111111111100000000000000000111110000011111110000001111111000000000000111111111111111", 
 "111111111111111100000000000000000111110000011111100000001111111000000000001111111111111111", 
 "111111111111111100001111000000000111110000011110000001111111100000000000011111111111111111", 
 "111111111111111100001111000000000111110000011110000001111111100000000000111111111111111111", 
 "111111111111111100001111000000000111100000011110000001111111100000000000111111111111111111", 
 "111111111111111100000011111111111110000000011110000111111111111111111000001111111111111111", 
 "111111111111111100000011111111111110000000011110000111111111111111111000000111111111111111", 
 "111111111111111100000010000000000000000000011110000001000000000000100000000111111111111111", 
 "111111111111111111100000000000000000000000011110000000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000011110000000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000011111000000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000001111111110000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000001111111110000000000000000000000001111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



fifty_three  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111000000000000000000000000000111111100000000000000000001111111111111111111111", 
 "111111111111111000000000000000000000000000111111100000000000000000001111111111111111111111", 
 "111111111111111000000000000000000000000000111111000000000000000000000111111111111111111111", 
 "111111111111111000000000000000000000000000111100000000000000000000000001111111111111111111", 
 "111111111111111000011111111111111111100000111100000011111111111110000001111111111111111111", 
 "111111111111111000011111000000000000000000111100000011100000001110000000011111111111111111", 
 "111111111111111000011110000000000000000000111100001111100000000111110000001111111111111111", 
 "111111111111111000011110000000000000000000111100001111000000000111110000001111111111111111", 
 "111111111111111000011111000000000000000000111100000000000000000111110000001111111111111111", 
 "111111111111111000011111111111111100000000111100000000000000000111110000001111111111111111", 
 "111111111111111000011111111111111100000000111100000000000000000111110000001111111111111111", 
 "111111111111111000000000000000001111100000111111100000000011111110000000011111111111111111", 
 "111111111111111000000000000000001111100000111111100000000011111110000000001111111111111111", 
 "111111111111111000000000000000001111100000111111000000000011111110000000001111111111111111", 
 "111111111111111000000000000000001111100000111100000000000000000111110000001111111111111111", 
 "111111111111111000000000000000001111100000111100000000000000000111110000001111111111111111", 
 "111111111111111000000000000000001111100000111100000000000000000111110000001111111111111111", 
 "111111111111111000011110000000001111100000111100001111100000000111110000001111111111111111", 
 "111111111111111000011110000000001111100000111100001111100000000111110000001111111111111111", 
 "111111111111111000000111111111111100000000111100000011111111111110000000011111111111111111", 
 "111111111111111000000111111111111100000000111100000011111111111110000000001111111111111111", 
 "111111111111111000000111111111111100000000111100000011111111111110000000001111111111111111", 
 "111111111111111111000000000000000000000000111111100000000000000000000000001111111111111111", 
 "111111111111111111000000000000000000000000111111100000000000000000000000001111111111111111", 
 "111111111111111111000000000000000000000000111111100000000000000000000000011111111111111111", 
 "111111111111111111111000000000000000000011111111111100000000000000000001111111111111111111", 
 "111111111111111111111000000000000000000011111111111100000000000000000001111111111111111111", 
 "111111111111111111111000000000000000000111111111111100000000000001000011111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



fifty_four   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111100000000000000000000000000011111111111111100000000000111111111111111111111", 
 "111111111111111100000000000000000000000000011111111111111100000000000111111111111111111111", 
 "111111111111111100000000000000000000000000011111111111111100000000000011111111111111111111", 
 "111111111111111100001111111111111111110000011111111111110000000000000000111111111111111111", 
 "111111111111111100001111111111111111100000011111111111110000011111000000111111111111111111", 
 "111111111111111100001111000000000000000000011111111111100000011111000000111111111111111111", 
 "111111111111111100001111000000000000000000011111111110000001111111000000111111111111111111", 
 "111111111111111100001111000000000000000000011111111110000001111111000000111111111111111111", 
 "111111111111111100001111111111111110000000011111110000000011111111000000111111111111111111", 
 "111111111111111100001111111111111110000000011111110000001111111111000000111111111111111111", 
 "111111111111111100000000000000001111000000011111110000001111111111000000111111111111111111", 
 "111111111111111100000000000000000111110000011110000001111100011111000000111111111111111111", 
 "111111111111111100000000000000000111110000011110000001111100011111000000111111111111111111", 
 "111111111111111100000000000000000111110000011110000001111100011111000000111111111111111111", 
 "111111111111111100000000000000000111110000011110000111110000011111000000111111111111111111", 
 "111111111111111100000000000000000111110000011110000111110000011111000000111111111111111111", 
 "111111111111111100001111000000000111110000011110000111110000011111000000001111111111111111", 
 "111111111111111100001111000000000111110000011110000111111111111111111000000111111111111111", 
 "111111111111111100000111000000000111000000011110000111111111111111111000000111111111111111", 
 "111111111111111100000011111111111110000000011110000000000000011111000000001111111111111111", 
 "111111111111111100000011111111111110000000011110000000000000011111000000000111111111111111", 
 "111111111111111100000000000000000000000000011110000000000000001111000000000111111111111111", 
 "111111111111111111100000000000000000000000011111100000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000011111110000000000000000000000000111111111111111", 
 "111111111111111111111000000000000000000000111111110000000000000000000000001111111111111111", 
 "111111111111111111111100000000000000000001111111111111111111000000000000111111111111111111", 
 "111111111111111111111100000000000000000001111111111111111111100000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



fifty_five   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111100000000000000000000000000011110000000000000000000000000000111111111111111", 
 "111111111111111100000000000000000000000000011110000000000000000000000000000111111111111111", 
 "111111111111111100000000000000000000000000011110000000000000000000000000000111111111111111", 
 "111111111111111100001111111111111111100000011110000111111111111111111000000111111111111111", 
 "111111111111111100001111111111111111110000011110000111111111111111111000000111111111111111", 
 "111111111111111100001111000000000000000000011110000111110000000000000000000111111111111111", 
 "111111111111111100001111000000000000000000011110000111110000000000000000000111111111111111", 
 "111111111111111100001111000000000000000000011110000111110000000000000000000111111111111111", 
 "111111111111111100001111111111111110000000011110000111111111111111000000000111111111111111", 
 "111111111111111100001111111111111110000000011110000111111111111111000000000111111111111111", 
 "111111111111111100000000000000001110000000011110000000000000000111000000001111111111111111", 
 "111111111111111100000000000000000111110000011110000000000000000011111000000111111111111111", 
 "111111111111111100000000000000000111110000011110000000000000000011111000000111111111111111", 
 "111111111111111100000000000000000111110000011110000000000000000011111000000111111111111111", 
 "111111111111111100000000000000000111110000011110000000000000000011111000000111111111111111", 
 "111111111111111100000000000000000111110000011110000000000000000011111000000111111111111111", 
 "111111111111111100001111000000000111110000011110000111100000000011111000000111111111111111", 
 "111111111111111100001111000000000111110000011110000111110000000011111000000111111111111111", 
 "111111111111111100001111000000000111100000011110000111110000000011110000001111111111111111", 
 "111111111111111100000011111111111110000000011110000001111111111111000000001111111111111111", 
 "111111111111111100000011111111111110000000011110000001111111111111000000000111111111111111", 
 "111111111111111100000000000000000000000000011110000000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000011111110000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000011111110000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000011111111000000000000000000000001111111111111111", 
 "111111111111111111111100000000000000000001111111111110000000000000000000111111111111111111", 
 "111111111111111111111100000000000000000001111111111110000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



fifty_six    <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111110000000000000000000000000001111111110000000000000111111111111111111111111", 
 "111111111111111110000000000000000000000000001111111110000000000000011111111111111111111111", 
 "111111111111111110000000000000000000000000001111111110000000000000011111111111111111111111", 
 "111111111111111110000111111111111111111000001111110000000000000000000011111111111111111111", 
 "111111111111111110000111111111111111110000001111110000001111111100000011111111111111111111", 
 "111111111111111110000111100000000000000000001111000000001110000000000011111111111111111111", 
 "111111111111111110000111100000000000000000001111000001111100000000000011111111111111111111", 
 "111111111111111110000111110000000000000000001110000001111100000000000011111111111111111111", 
 "111111111111111110000111111111111111000000001110000001110000000000000011111111111111111111", 
 "111111111111111110000111111111111111000000001110000111110000000000000011111111111111111111", 
 "111111111111111110000000000000000011110000001111000111110000000000000011111111111111111111", 
 "111111111111111110000000000000000011111000001111000111111111111111000000111111111111111111", 
 "111111111111111110000000000000000011111000001110000111111111111111000000011111111111111111", 
 "111111111111111110000000000000000011111000001110000111110000000111000000001111111111111111", 
 "111111111111111110000000000000000011111000001110000111110000000011111000000111111111111111", 
 "111111111111111110000000000000000011111000001110000111110000000011111000000111111111111111", 
 "111111111111111110000111100000000011111000001110000111110000000011111000000111111111111111", 
 "111111111111111110000111100000000011111000001110000111110000000011111000000111111111111111", 
 "111111111111111110000001111111111111000000001110000111110000000011111000000111111111111111", 
 "111111111111111110000001111111111111000000001111000001111111111111000000000111111111111111", 
 "111111111111111110000001111111111111000000001110000001111111111111000000000111111111111111", 
 "111111111111111111000000000000000000000000001111000001111111111111000000000111111111111111", 
 "111111111111111111110000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000000111111111000000000000000000000000111111111111111", 
 "111111111111111111111110000000000000000000111111111110000000000000000000011111111111111111", 
 "111111111111111111111110000000000000000000111111111110000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111000111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



fifty_seven  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111000001000000000000100000001111111111111111111111111111111111111111111111", 
 "111111111111111110000000000000000000000000001111100000000000000000000000011111111111111111", 
 "111111111111111110000000000000000000000000001111000000000000000000000000011111111111111111", 
 "111111111111111110000000000000000000000000001111000000000000000000000000001111111111111111", 
 "111111111111111110000111111111111111111000001111000000000000000000010000000111111111111111", 
 "111111111111111110000111111111111111110000001111000011111111111111111100000011111111111111", 
 "111111111111111110000111100000000000000000001111000011111111111111111000000011111111111111", 
 "111111111111111110000111100000000000000000001111000000000000001111100000000011111111111111", 
 "111111111111111110000111110000000000000000001111000000000000001111100000000011111111111111", 
 "111111111111111110000111111111111111000000001111100000000000001111100000000011111111111111", 
 "111111111111111110000111111111111111000000001111111000000000001111100000000011111111111111", 
 "111111111111111110000000000000000011100000001111111000000000001111100000000111111111111111", 
 "111111111111111110000000000000000011111000001111111111110000111100000000001111111111111111", 
 "111111111111111110000000000000000011111000001111111111111000111100000000011111111111111111", 
 "111111111111111110000000000000000011111000001111111111111000111100000000011111111111111111", 
 "111111111111111110000000000000000011111000001111111111000000111100000000011111111111111111", 
 "111111111111111110000000000000000011111000001111111111000000111100000000011111111111111111", 
 "111111111111111110000111100000000011111000001111111111000001110000000000011111111111111111", 
 "111111111111111110000111100000000011111000001111111111000111110000000011111111111111111111", 
 "111111111111111110000001110000000111000000001111111111000111110000000011111111111111111111", 
 "111111111111111110000001111111111111000000001111111111000111110000000011111111111111111111", 
 "111111111111111110000001111111111111000000001111111111000111110000000011111111111111111111", 
 "111111111111111110000000000000000000000000001111111111000000000000000011111111111111111111", 
 "111111111111111111110000000000000000000000001111111111000000000000011111111111111111111111", 
 "111111111111111111110000000000000000000000001111111111000000000000011111111111111111111111", 
 "111111111111111111111100000000000000000000111111111111000000000000011111111111111111111111", 
 "111111111111111111111110000000000000000000111111111111111000000000011111111111111111111111", 
 "111111111111111111111110000000000000000000111111111111111000000000011111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




fifty_eight  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111000001000000000000100000001111111001000000000000100111111111111111111111", 
 "111111111111111110000000000000000000000000001111110000000000000000000011111111111111111111", 
 "111111111111111110000000000000000000000000001111110000000000000000000011111111111111111111", 
 "111111111111111110000000000000000000000000001111000000000000000000000000111111111111111111", 
 "111111111111111110000111111111111111111000001111000001111111111111000000011111111111111111", 
 "111111111111111110000111111111111111111000001110000011110000000011111000000111111111111111", 
 "111111111111111110000111100000000000000000001110000111110000000011111000000111111111111111", 
 "111111111111111110000111100000000000000000001110000111110000000011111000000111111111111111", 
 "111111111111111110000111110000000000000000001110000111110000000011111000000111111111111111", 
 "111111111111111110000111111111111111000000001110000111111100000011111000000111111111111111", 
 "111111111111111110000111111111111111000000001111000111111100000011111000000111111111111111", 
 "111111111111111110000000000000000011100000001111000001111110000011100000000111111111111111", 
 "111111111111111110000000000000000011111000001111000001111111111111000000000111111111111111", 
 "111111111111111110000000000000000011111000001110000001111111111111000000000111111111111111", 
 "111111111111111110000000000000000011111000001110000011110000011111110000000111111111111111", 
 "111111111111111110000000000000000011111000001110000111110000001111111000000111111111111111", 
 "111111111111111110000000000000000011111000001110000111110000000011111000000111111111111111", 
 "111111111111111110000111100000000011111000001110000111110000000011111000000111111111111111", 
 "111111111111111110000111100000000011111000001110000111110000000011111000000111111111111111", 
 "111111111111111110000001110000000111000000001111000001110000000011100000000111111111111111", 
 "111111111111111110000001111111111111000000001111000001111111111111000000000111111111111111", 
 "111111111111111110000001111111111111000000001110000001111111111111000000000111111111111111", 
 "111111111111111110000000000000000000000000001111000000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000000111111111110000000000000000000011111111111111111", 
 "111111111111111111111110000000000000000000111111111110000000000000000000011111111111111111", 
 "111111111111111111111110000000000000000000111111111110000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




fifty_nine   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111100000000000000000000000000011111110000000000000000000111111111111111111111", 
 "111111111111111100000000000000000000000000011111110000000000000000000111111111111111111111", 
 "111111111111111100000000000000000000000000011111100000000000000000000011111111111111111111", 
 "111111111111111100000010000000000001000000011110000000000000000000000000111111111111111111", 
 "111111111111111100001111111111111111110000011110000001111111111111000000111111111111111111", 
 "111111111111111100001111100000000000000000011110000001110000000011000000001111111111111111", 
 "111111111111111100001111000000000000000000011110000111110000000011111000000111111111111111", 
 "111111111111111100001111000000000000000000011110000111110000000011111000000111111111111111", 
 "111111111111111100001111111111111100000000011110000111110000000011111000000111111111111111", 
 "111111111111111100001111111111111110000000011110000111110000000011111000000111111111111111", 
 "111111111111111100001111111111111110000000011110000111110000000011111000000111111111111111", 
 "111111111111111100000000000000000111110000011110000001111111111111111000001111111111111111", 
 "111111111111111100000000000000000111110000011110000001111111111111111000000111111111111111", 
 "111111111111111100000000000000000111110000011110000001111111111111111000000111111111111111", 
 "111111111111111100000000000000000111110000011111110000000000000011111000000111111111111111", 
 "111111111111111100000000000000000111110000011111110000000000000011111000000111111111111111", 
 "111111111111111100000000000000000111110000011111111000000000000111000000000111111111111111", 
 "111111111111111100001111000000000111110000011111111110000000011111000000000111111111111111", 
 "111111111111111100001111000000000111100000011111111110000000011111000000000111111111111111", 
 "111111111111111100000011111111111110000000011111111110001111111000000000001111111111111111", 
 "111111111111111100000011111111111110000000011111111110001111111000000000000111111111111111", 
 "111111111111111100000011111111111110000000011111111110001111111000000000000111111111111111", 
 "111111111111111111100000000000000000000000011111111110000000000000000000111111111111111111", 
 "111111111111111111100000000000000000000000011111111110000000000000000000111111111111111111", 
 "111111111111111111100000000000000000000000011111111110000000000000000000111111111111111111", 
 "111111111111111111111100000000000000000001111111111111110000000000000111111111111111111111", 
 "111111111111111111111100000000000000000001111111111111110000000000000111111111111111111111", 
 "111111111111111111111110000000000011000011111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




sixty        <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111000000000000000000111111111111111111111", 
 "111111111111111111111000000000000011111111111111110000000000000000000111111111111111111111", 
 "111111111111111111111000000000000011111111111111100000000000000000000111111111111111111111", 
 "111111111111111111100000000000000000011111111110000000000000000000000000111111111111111111", 
 "111111111111111111000000111111100000001111111110000001111111111111000000111111111111111111", 
 "111111111111111111000000111111100000001111111110000001110000000111000000001111111111111111", 
 "111111111111111100000000110000000000001111111110000111100000000011111000000111111111111111", 
 "111111111111111000000111110000000000001111111110000111100000000011111000000111111111111111", 
 "111111111111111000000111110000000000001111111110000111100000000111111000000111111111111111", 
 "111111111111111000011111000000000000001111111110000111100000011111111000000111111111111111", 
 "111111111111111000011111000000000000001111111110000111100000011111111000000111111111111111", 
 "111111111111111000011111000000000000001111111111000111110001100011111000000111111111111111", 
 "111111111111111000011111111111111100000011111110000111100001100011111000000111111111111111", 
 "111111111111111000011111111111111100000011111110000111110001000011111000000111111111111111", 
 "111111111111111000011111000000001100000000111110000111111100000011111000000111111111111111", 
 "111111111111111000011111000000001111100000011110000111111100000011111000000111111111111111", 
 "111111111111111000011111000000001111100000011110000111110000000011111000000111111111111111", 
 "111111111111111000011111000000001111100000011110000111100000000011111000000111111111111111", 
 "111111111111111000011111000000001111100000011110000111100000000011111000000111111111111111", 
 "111111111111111000011111000000001111100000011111000001111111111111000000000111111111111111", 
 "111111111111111000000111111111111100000000011110000001111111111111000000000111111111111111", 
 "111111111111111000000111111111111100000000011110000001111111111111000000000111111111111111", 
 "111111111111111000000111111111111100000000011111110000000000000000000000000111111111111111", 
 "111111111111111111000000000000000000000000011111110000000000000000000000000111111111111111", 
 "111111111111111111000000000000000000000000011111110000000000000000000000001111111111111111", 
 "111111111111111111100000000000000000000000111111111100000000000000000000111111111111111111", 
 "111111111111111111111000000000000000000011111111111110000000000000000000111111111111111111", 
 "111111111111111111111000000000000010000011111111111110000000000000000001111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");





sixty_one    <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111100000000000111111111111111111111111", 
 "111111111111111111111100000000000001111111111111111111100000000000111111111111111111111111", 
 "111111111111111111111100000000000001111111111111111110000000000000001111111111111111111111", 
 "111111111111111111100000000000000000001111111111111100000011111000000111111111111111111111", 
 "111111111111111111100000011111110000000111111111111100000011111000000111111111111111111111", 
 "111111111111111111100000011111110000000111111111111100000011111000000111111111111111111111", 
 "111111111111111100000011111000000000000111111111111100011111111000000111111111111111111111", 
 "111111111111111100000011111000000000000111111111111100000011111000000111111111111111111111", 
 "111111111111111100000011100000000000000111111111111100000011111000000111111111111111111111", 
 "111111111111111100001111100000000000000111111111111100000011111000000111111111111111111111", 
 "111111111111111100001111100000000000000111111111111110000011111000000111111111111111111111", 
 "111111111111111100001111111111111110000001111111111111100011111000000111111111111111111111", 
 "111111111111111100001111111111111110000001111111111111100011111000000111111111111111111111", 
 "111111111111111100001111111111111110000001111111111111100011111000000111111111111111111111", 
 "111111111111111100001111100000000111100000001111111111100011111000000111111111111111111111", 
 "111111111111111100001111100000000111110000001111111111100011111000000111111111111111111111", 
 "111111111111111100001111100000000111110000001111110000000011111000000000111111111111111111", 
 "111111111111111100001111100000000111110000001111110000000011111000000000111111111111111111", 
 "111111111111111100001111100000000111110000001111110000000011111000000000111111111111111111", 
 "111111111111111100000011100000000111000000001111110001111111111111111000000111111111111111", 
 "111111111111111100000011111111111110000000001111110001111111111111110000000111111111111111", 
 "111111111111111100000011111111111110000000001111110000000000000000000000000111111111111111", 
 "111111111111111110000000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000001111111000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000000111111111100000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000001111111111100000000000000000000000111111111111111", 
 "111111111111111111111100000111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");





sixty_two    <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111110000000000000000000111111111111111111111", 
 "111111111111111111111100000000000001111111111111110000000000000000000011111111111111111111", 
 "111111111111111111111100000000000001111111111111000000000000000000000000111111111111111111", 
 "111111111111111111100000000000000000001111111111000000111111111111000000111111111111111111", 
 "111111111111111111100000011111110000000111111111000001111111111111000000011111111111111111", 
 "111111111111111111100000011111110000000111111111000001110000000011100000000111111111111111", 
 "111111111111111100000011111000000000000111111111000111110000000011111000000111111111111111", 
 "111111111111111100000011111000000000000111111111000111110000000011111000000111111111111111", 
 "111111111111111100000011100000000000000111111111000111110000001111111000000111111111111111", 
 "111111111111111100001111100000000000000111111111000111110000001111111000000111111111111111", 
 "111111111111111100001111100000000000000111111111000111100000011111111000000111111111111111", 
 "111111111111111100001111100000000000000001111111000000000001111111000000000111111111111111", 
 "111111111111111100001111111111111110000001111111000000000001111111000000000111111111111111", 
 "111111111111111100001111111111111110000001111111000000000001111100000000000111111111111111", 
 "111111111111111100001111100000000111000000011111110000001111111100000000000111111111111111", 
 "111111111111111100001111100000000111110000001111110000001111111000000000000111111111111111", 
 "111111111111111100001111100000000111110000001111000000111111100000000000011111111111111111", 
 "111111111111111100001111100000000111110000001111000001111111100000000000011111111111111111", 
 "111111111111111100001111100000000111110000001111000001111111100000000000011111111111111111", 
 "111111111111111100000011100000000111000000001111000111111111111111111000000111111111111111", 
 "111111111111111100000011111111111110000000001111000111111111111111111000000111111111111111", 
 "111111111111111100000011111111111110000000001111000001000000000000100000000111111111111111", 
 "111111111111111110000000000000000000000000001111000000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000001111000000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000001111000000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000000111111110000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000001111111110000000000000000000000000111111111111111", 
 "111111111111111111111100000111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");





sixty_three  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111110000000000000111111111111111100000000000000000011111111111111111111", 
 "111111111111111111111110000000000000111111111111111000000000000000000001111111111111111111", 
 "111111111111111111111110000000000000011111111111111000000000000000000001111111111111111111", 
 "111111111111111111110000000000000000000111111111100000000000000000000000011111111111111111", 
 "111111111111111111110000001111111000000011111111100000111111111111100000001111111111111111", 
 "111111111111111111000000001110000000000011111111100000111000000001100000000111111111111111", 
 "111111111111111110000001111100000000000011111111100011111000000001111100000011111111111111", 
 "111111111111111110000001111100000000000011111111100011111000000001111100000011111111111111", 
 "111111111111111110000001110000000000000011111111100000000000000001111100000011111111111111", 
 "111111111111111110000111110000000000000011111111100000000000000001111100000011111111111111", 
 "111111111111111110000111110000000000000011111111100000000000000001111100000011111111111111", 
 "111111111111111110000111111111111111000000111111111000000000111111100000000011111111111111", 
 "111111111111111110000111111111111111000000111111111000000000111111100000000011111111111111", 
 "111111111111111110000111111111111111000000011111111000000000111111100000000011111111111111", 
 "111111111111111110000111110000000011111000000111100000000000000001111100000011111111111111", 
 "111111111111111110000111110000000011111000000111100000000000000001111100000011111111111111", 
 "111111111111111110000111110000000011111000000111100000000000000001111100000011111111111111", 
 "111111111111111110000111110000000011111000000111100011111000000001111100000011111111111111", 
 "111111111111111110000111110000000011111000000111100011111000000001111100000011111111111111", 
 "111111111111111110000001111111111111000000000111100000111111111111110000000011111111111111", 
 "111111111111111110000001111111111111000000000111100000111111111111100000000011111111111111", 
 "111111111111111110000001111111111111000000000111100000111111111111100000000011111111111111", 
 "111111111111111111110000000000000000000000000111111000000000000000000000000011111111111111", 
 "111111111111111111110000000000000000000000000111111000000000000000000000000011111111111111", 
 "111111111111111111110000000000000000000000001111111100000000000000000000000011111111111111", 
 "111111111111111111111110000000000000000000111111111111000000000000000000001111111111111111", 
 "111111111111111111111110000000000000000000111111111111000000000000000000011111111111111111", 
 "111111111111111111111111000111111111111111111111111111100000000000000000011111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");





sixty_four   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111110000000000111111111111111111111", 
 "111111111111111111111100000000000001111111111111111111111100000000000011111111111111111111", 
 "111111111111111111111100000000000001111111111111111111111100000000000011111111111111111111", 
 "111111111111111111110000000000000000001111111111111111110000000000000000111111111111111111", 
 "111111111111111111100000011111110000000111111111111111110000001111000000011111111111111111", 
 "111111111111111111100000011111110000000111111111111111110000011111000000011111111111111111", 
 "111111111111111110000000011100000000000111111111111110000001111111000000011111111111111111", 
 "111111111111111100000011111000000000000111111111111110000001111111000000011111111111111111", 
 "111111111111111100000011110000000000000111111111110000000011111111000000011111111111111111", 
 "111111111111111100001111100000000000000111111111110000001111111111000000011111111111111111", 
 "111111111111111100001111100000000000000111111111110000001111111111000000111111111111111111", 
 "111111111111111100001111100000000000000011111111000000111110011111000000111111111111111111", 
 "111111111111111100001111111111111110000001111111000001111100001111000000011111111111111111", 
 "111111111111111100001111111111111110000001111111000001111100001111000000011111111111111111", 
 "111111111111111100001111100000000110000000011111000111110000001111000000011111111111111111", 
 "111111111111111100001111100000000111110000001111000111110000001111000000011111111111111111", 
 "111111111111111100001111100000000111110000001111000111110000011111100000000111111111111111", 
 "111111111111111100001111100000000111110000001111000111111111111111111000000111111111111111", 
 "111111111111111100001111100000000111110000001111000111111111111111111000000111111111111111", 
 "111111111111111100001111100000000111110000001111000000000000011111100000000111111111111111", 
 "111111111111111100000011111111111110000000001111000000000000001111000000000111111111111111", 
 "111111111111111100000011111111111110000000001111000000000000001111000000000111111111111111", 
 "111111111111111100000000000000000000000000001111100000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000001111111000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000011111111111111111100000000000011111111111111111", 
 "111111111111111111111100000000000000000001111111111111111111100000000000011111111111111111", 
 "111111111111111111111100000111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");





sixty_five   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111000000000000111111111111100000000000000000000000000011111111111111", 
 "111111111111111111111110000000000000111111111111100000000000000000000000000011111111111111", 
 "111111111111111111111110000000000000011111111111100000000000000000000000000011111111111111", 
 "111111111111111111110000000000000000000111111111100011111111111111111100000011111111111111", 
 "111111111111111111110000001111111000000011111111100011111111111111111100000011111111111111", 
 "111111111111111111000000001110000000000011111111100011111000000000000000000011111111111111", 
 "111111111111111110000001111100000000000011111111100011111000000000000000000011111111111111", 
 "111111111111111110000001111100000000000011111111100011111000000000000000000011111111111111", 
 "111111111111111110000001110000000000000011111111100011111111111111100000000011111111111111", 
 "111111111111111110000111110000000000000011111111100011111111111111100000000011111111111111", 
 "111111111111111110000111110000000000000011111111100000000000000011110000000011111111111111", 
 "111111111111111111000111111111111111000000111111100000000000000001111100000011111111111111", 
 "111111111111111110000111111111111111000000111111100000000000000001111100000011111111111111", 
 "111111111111111110000111111111111111000000011111100000000000000001111100000011111111111111", 
 "111111111111111110000111110000000011111000000111100000000000000001111100000011111111111111", 
 "111111111111111110000111110000000011111000000111100000000000000001111100000011111111111111", 
 "111111111111111110000111110000000011111000000111100011111000000001111100000011111111111111", 
 "111111111111111110000111110000000011111000000111100011111000000001111100000011111111111111", 
 "111111111111111110000111110000000011111000000111100011111000000001111100000011111111111111", 
 "111111111111111110000001111111111111000000000111100000111111111111100000000011111111111111", 
 "111111111111111110000001111111111111000000000111100000111111111111100000000011111111111111", 
 "111111111111111110000001111111111111000000000111100000000000000000000000000011111111111111", 
 "111111111111111111110000000000000000000000000111111000000000000000000000000011111111111111", 
 "111111111111111111110000000000000000000000000111111000000000000000000000000011111111111111", 
 "111111111111111111110000000000000000000000001111111100000000000000000000000111111111111111", 
 "111111111111111111111110000000000000000000111111111111000000000000000000001111111111111111", 
 "111111111111111111111110000000000000000000111111111111000000000000000000011111111111111111", 
 "111111111111111111111110000111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");





sixty_six    <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111000000000000011111111111111111100000000000001111111111111111111111", 
 "111111111111111111111111000000000000011111111111111111000000000000001111111111111111111111", 
 "111111111111111111111110000000000000001111111111111111000000000000001111111111111111111111", 
 "111111111111111111111000000000000000000001111111111000000000000000000001111111111111111111", 
 "111111111111111111111000000111111100000001111111111000000111111110000001111111111111111111", 
 "111111111111111111100000000111000000000001111111100000000111000000000001111111111111111111", 
 "111111111111111111000000111110000000000001111111100000011111000000000001111111111111111111", 
 "111111111111111111000000111110000000000001111111100000011111000000000001111111111111111111", 
 "111111111111111111000001111000000000000001111111100000111000000000000001111111111111111111", 
 "111111111111111111000011111000000000000001111111100011111000000000000001111111111111111111", 
 "111111111111111111000011111000000000000001111111100011111000000000000001111111111111111111", 
 "111111111111111111000011111111111111100000011111100011111111111111110000001111111111111111", 
 "111111111111111111000011111111111111100000011111100011111111111111100000001111111111111111", 
 "111111111111111111000011111000000011100000000111100011111100000001110000000111111111111111", 
 "111111111111111111000011111000000001111100000011100011111000000000111100000011111111111111", 
 "111111111111111111000011111000000001111100000011100011111000000000111100000011111111111111", 
 "111111111111111111000011111000000001111100000011100011111000000000111100000011111111111111", 
 "111111111111111111000011111000000001111100000011100011111000000000111100000011111111111111", 
 "111111111111111111000011111000000001111100000011100011111000000000111100000011111111111111", 
 "111111111111111111000000111111111111100000000111100000011111111111110000000011111111111111", 
 "111111111111111111000000111111111111100000000011100000011111111111100000000011111111111111", 
 "111111111111111111000000111111111111100000000011100000011111111111100000000011111111111111", 
 "111111111111111111111000000000000000000000000011111000000000000000000000000011111111111111", 
 "111111111111111111111000000000000000000000000011111000000000000000000000000011111111111111", 
 "111111111111111111111000000000000000000000000111111100000000000000000000000011111111111111", 
 "111111111111111111111111000000000000000000011111111111000000000000000000001111111111111111", 
 "111111111111111111111111000000000000000000011111111111000000000000000000011111111111111111", 
 "111111111111111111111111100011111111111111111111111111100011111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");





sixty_seven  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111100000000000001111111111111000000000000000000000000111111111111111111", 
 "111111111111111111111100000000000001111111111111000000000000000000000000011111111111111111", 
 "111111111111111111111100000000000000111111111111000000000000000000000000011111111111111111", 
 "111111111111111111100000000000000000001111111111000000000000000000000000000111111111111111", 
 "111111111111111111100000011111110000000111111111000111111111111111111000000111111111111111", 
 "111111111111111111100000011111110000000111111111000111111111111111111000000111111111111111", 
 "111111111111111100000011111000000000000111111111000000000000001111000000000111111111111111", 
 "111111111111111100000011111000000000000111111111000000000000001111000000000111111111111111", 
 "111111111111111100000011100000000000000111111111000000000000001111000000000111111111111111", 
 "111111111111111100001111100000000000000111111111110000000000001111000000000111111111111111", 
 "111111111111111100001111100000000000000111111111110000000000011111000000000111111111111111", 
 "111111111111111100001111111111111110000001111111111111110001111100000000011111111111111111", 
 "111111111111111100001111111111111110000001111111111111110001111100000000111111111111111111", 
 "111111111111111100001111111111111110000000111111111111110001111100000000011111111111111111", 
 "111111111111111100001111100000000111110000001111111110000001111100000000011111111111111111", 
 "111111111111111100001111100000000111110000001111111110000001111000000000011111111111111111", 
 "111111111111111100001111100000000111110000001111111110000001100000000000111111111111111111", 
 "111111111111111100001111100000000111110000001111111110001111100000000011111111111111111111", 
 "111111111111111100001111100000000111110000001111111110001111100000000111111111111111111111", 
 "111111111111111100000011111111111110000000001111111110001111100000000011111111111111111111", 
 "111111111111111100000011111111111110000000001111111110001111100000000011111111111111111111", 
 "111111111111111100000011111111111110000000001111111110000000000000000111111111111111111111", 
 "111111111111111111000000000000000000000000001111111110000000000000011111111111111111111111", 
 "111111111111111111100000000000000000000000001111111110000000000000011111111111111111111111", 
 "111111111111111111100000000000000000000000011111111110000000000000011111111111111111111111", 
 "111111111111111111111100000000000000000001111111111111110000000000011111111111111111111111", 
 "111111111111111111111100000000000000000001111111111111110000000000011111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");





sixty_eight  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111100000000000001111111111111110010000000000001001111111111111111111111", 
 "111111111111111111111100000000000001111111111111100000000000000000000111111111111111111111", 
 "111111111111111111100000000000000000001111111111100000000000000000000111111111111111111111", 
 "111111111111111111100000011111110000000111111110000000000000000000000000111111111111111111", 
 "111111111111111111100000011111110000000111111110000001111111111110000000111111111111111111", 
 "111111111111111100000011111000000000000111111110000111100000000111110000001111111111111111", 
 "111111111111111100000011111000000000000111111110001111100000000011110000001111111111111111", 
 "111111111111111100000011100000000000000111111110001111100000000011110000001111111111111111", 
 "111111111111111100001111100000000000000111111110001111110000000011110000001111111111111111", 
 "111111111111111100001111100000000000000111111110001111111100000011110000001111111111111111", 
 "111111111111111100001111100000000000000011111110001111111100000011110000001111111111111111", 
 "111111111111111100001111111111111110000001111110000011111100000111000000001111111111111111", 
 "111111111111111100001111111111111110000001111110000001111111111110000000001111111111111111", 
 "111111111111111100001111100000000111000000011110000001111111111110000000001111111111111111", 
 "111111111111111100001111100000000111110000001110000111100000011111110000001111111111111111", 
 "111111111111111100001111100000000111110000001110001111100000011111110000001111111111111111", 
 "111111111111111100001111100000000111110000001110001111100000000111110000001111111111111111", 
 "111111111111111100001111100000000111110000001110001111100000000011110000001111111111111111", 
 "111111111111111100001111100000000111100000001110001111100000000011110000001111111111111111", 
 "111111111111111100000011111111111110000000001110000011100000000111000000001111111111111111", 
 "111111111111111100000011111111111110000000001110000001111111111110000000001111111111111111", 
 "111111111111111110000000000000000000000000001110000001111111111110000000001111111111111111", 
 "111111111111111111100000000000000000000000001110000000000000000000000000001111111111111111", 
 "111111111111111111100000000000000000000000001111100000000000000000000000001111111111111111", 
 "111111111111111111110000000000000000000000011111110000000000000000000000001111111111111111", 
 "111111111111111111111100000000000000000001111111111100000000000000000000111111111111111111", 
 "111111111111111111111100000111111111111111111111111100000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111110000000000000000001111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");





sixty_nine   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111110000000000000111111111111111000000000000000000011111111111111111111", 
 "111111111111111111111110000000000000111111111111111000000000000000000001111111111111111111", 
 "111111111111111111111100000000000000011111111111110000000000000000000001111111111111111111", 
 "111111111111111111110000000000000000000011111111100000000000000000000000011111111111111111", 
 "111111111111111111110000001111111000000011111111100000111111111111100000001111111111111111", 
 "111111111111111111000000001110000000000011111111100000111000000001110000000011111111111111", 
 "111111111111111110000001111100000000000011111111100011111000000001111100000011111111111111", 
 "111111111111111110000001111100000000000011111111100011111000000001111100000011111111111111", 
 "111111111111111110000011110000000000000011111111100011111000000001111100000011111111111111", 
 "111111111111111110000111110000000000000011111111100011111000000001111100000011111111111111", 
 "111111111111111110000111110000000000000011111111100011111000000001111100000011111111111111", 
 "111111111111111110000111111111111111000000111111100000111111111111111100000011111111111111", 
 "111111111111111110000111111111111111000000111111100000111111111111111100000011111111111111", 
 "111111111111111110000111111111111111000000011111100000011111111111111100000011111111111111", 
 "111111111111111110000111110000000011111000000111111000000000000001111100000011111111111111", 
 "111111111111111110000111110000000011111000000111111000000000000001111100000011111111111111", 
 "111111111111111110000111110000000011111000000111111100000000000001100000000011111111111111", 
 "111111111111111110000111110000000011111000000111111111000000000111100000000011111111111111", 
 "111111111111111110000111110000000011111000000111111111000000001111100000000011111111111111", 
 "111111111111111110000001111111111111000000000111111111000111111110000000000011111111111111", 
 "111111111111111110000001111111111111000000000111111111000111111110000000000011111111111111", 
 "111111111111111110000001111111111111000000000111111111000111111100000000000011111111111111", 
 "111111111111111111110000000000000000000000000111111111000000000000000000001111111111111111", 
 "111111111111111111110000000000000000000000000111111111000000000000000000011111111111111111", 
 "111111111111111111110000000000000000000000001111111111000000000000000000011111111111111111", 
 "111111111111111111111110000000000000000000111111111111111000000000000001111111111111111111", 
 "111111111111111111111110000000000000000000111111111111111000000000000011111111111111111111", 
 "111111111111111111111111101111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");





seventy      <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111110000000000000000000000001111111111000000000000000000111111111111111111111", 
 "111111111111111100000000000000000000000001111111110000000000000000000011111111111111111111", 
 "111111111111111100000000000000000000000000111111110000000000000000000011111111111111111111", 
 "111111111111111100000010000000000000000000001111000000000000000000000000111111111111111111", 
 "111111111111111100001111111111111111110000001111000001111111111111000000011111111111111111", 
 "111111111111111100000010000000111111000000001111000001110000000111000000001111111111111111", 
 "111111111111111100000000000000111110000000001111000111110000000011111000000111111111111111", 
 "111111111111111100000000000000111110000000001111000111110000000011111000000111111111111111", 
 "111111111111111110000000000000111110000000001111000111110000000011111000000111111111111111", 
 "111111111111111111100000000000111110000000001111000111110000001111111000000111111111111111", 
 "111111111111111111100000000000111110000000001111000111110000001111111000000111111111111111", 
 "111111111111111111111111100011111000000001111111000111110001100011111000000111111111111111", 
 "111111111111111111111111100011110000000001111111000111110001100011111000000111111111111111", 
 "111111111111111111111111000011110000000001111111000111110000100011111000000111111111111111", 
 "111111111111111111111100000011110000000001111111000111111100000011111000000111111111111111", 
 "111111111111111111111100000011110000000001111111000111111100000011111000000111111111111111", 
 "111111111111111111111100000011000000000001111111000111110000000011111000000111111111111111", 
 "111111111111111111111100011111000000000111111111000111110000000011111000000111111111111111", 
 "111111111111111111111100011111000000000111111111000111110000000011111000000111111111111111", 
 "111111111111111111111100011111000000000111111111000001111111111111100000000111111111111111", 
 "111111111111111111111100011111000000000111111111000001111111111111000000000111111111111111", 
 "111111111111111111111100000000000000001111111111000001111111111111000000000111111111111111", 
 "111111111111111111111100000000000000111111111111110000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000111111111111110000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000111111111111110000000000000000000000000111111111111111", 
 "111111111111111111111111000000000000111111111111111110000000000000000000011111111111111111", 
 "111111111111111111111111100000000000111111111111111110000000000000000000011111111111111111", 
 "111111111111111111111111100000000001111111111111111111000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




seventy_one  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111100000000000000000000000001111111111111000000000000111111111111111111111111", 
 "111111111111111100000000000000000000000001111111111111000000000000111111111111111111111111", 
 "111111111111111100000000000000000000000000011111111100000000000000001111111111111111111111", 
 "111111111111111100001111111111111111110000001111111100000011110000001111111111111111111111", 
 "111111111111111100001111111111111111110000001111111100000011110000001111111111111111111111", 
 "111111111111111100000000000000111110000000001111111100000011110000001111111111111111111111", 
 "111111111111111100000000000000111110000000001111111100011111110000001111111111111111111111", 
 "111111111111111100000000000000111110000000001111111100000111110000001111111111111111111111", 
 "111111111111111111100000000000111110000000001111111100000011110000001111111111111111111111", 
 "111111111111111111100000000000111110000000001111111100000011110000001111111111111111111111", 
 "111111111111111111110000000000111000000000011111111100000011110000001111111111111111111111", 
 "111111111111111111111111100011110000000001111111111111000011110000001111111111111111111111", 
 "111111111111111111111111100011110000000001111111111111000011110000001111111111111111111111", 
 "111111111111111111111100000011110000000001111111111111000011110000001111111111111111111111", 
 "111111111111111111111100000011110000000001111111111111000011110000001111111111111111111111", 
 "111111111111111111111100000011110000000001111111111111000011110000001111111111111111111111", 
 "111111111111111111111100001111000000000111111111100000000011110000000001111111111111111111", 
 "111111111111111111111100011111000000000111111111100000000011110000000001111111111111111111", 
 "111111111111111111111100011111000000000111111111100000000011111000000001111111111111111111", 
 "111111111111111111111100011111000000000111111111100011111111111111110000001111111111111111", 
 "111111111111111111111100001111000000000111111111100011111111111111110000001111111111111111", 
 "111111111111111111111100000000000000111111111111100000000000000000000000001111111111111111", 
 "111111111111111111111100000000000000111111111111100000000000000000000000001111111111111111", 
 "111111111111111111111100000000000000111111111111100000000000000000000000001111111111111111", 
 "111111111111111111111110000000000000111111111111110000000000000000000000001111111111111111", 
 "111111111111111111111111100000000000111111111111111100000000000000000000001111111111111111", 
 "111111111111111111111111100000000000111111111111111100000000000000000000001111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




seventy_two  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111110000000000000000000000001111111110000000000000000000111111111111111111111", 
 "111111111111111100000000000000000000000001111111100000000000000000000111111111111111111111", 
 "111111111111111100000000000000000000000000011110000000000000000000000001111111111111111111", 
 "111111111111111100001111111111111111110000001110000001111111111110000000111111111111111111", 
 "111111111111111100001111111111111111110000001110000001111111111111000000111111111111111111", 
 "111111111111111100000000000000111110000000001110000011100000000111000000001111111111111111", 
 "111111111111111100000000000000111110000000001110001111100000000011111000001111111111111111", 
 "111111111111111100000000000000111110000000001110001111100000000111111000001111111111111111", 
 "111111111111111111100000000000111110000000001110001111100000011111111000001111111111111111", 
 "111111111111111111100000000000111110000000001110001111100000011111111000001111111111111111", 
 "111111111111111111100000000000111100000000001110000111100000011111110000001111111111111111", 
 "111111111111111111111111100011111000000001111110000000000011111111000000001111111111111111", 
 "111111111111111111111111100011110000000001111110000000000011111111000000001111111111111111", 
 "111111111111111111111100000011110000000001111110000000000011111000000000001111111111111111", 
 "111111111111111111111100000011110000000001111111100000001111111000000000001111111111111111", 
 "111111111111111111111100000011110000000001111111100000011111110000000000001111111111111111", 
 "111111111111111111111100001111000000000111111110000001111111000000000000111111111111111111", 
 "111111111111111111111100011111000000000111111110000001111111000000000000111111111111111111", 
 "111111111111111111111100011111000000001111111110000001111111000000000000111111111111111111", 
 "111111111111111111111100011111000000000111111110001111111111111111111000001111111111111111", 
 "111111111111111111111100011111000000000111111110001111111111111111111000001111111111111111", 
 "111111111111111111111100000000000000111111111110000010000000000001100000001111111111111111", 
 "111111111111111111111100000000000000111111111110000000000000000000000000001111111111111111", 
 "111111111111111111111100000000000000111111111110000000000000000000000000001111111111111111", 
 "111111111111111111111110000000000000111111111111000000000000000000000000001111111111111111", 
 "111111111111111111111111100000000000111111111111100000000000000000000000001111111111111111", 
 "111111111111111111111111100000000000111111111111110000000000000000000000001111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




seventy_three<=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111110000000000000000000000001111111110000000000000000000111111111111111111111", 
 "111111111111111100000000000000000000000001111111100000000000000000000111111111111111111111", 
 "111111111111111100000000000000000000000000111111100000000000000000000111111111111111111111", 
 "111111111111111100000010000000000000000000001110000000000000000000000000111111111111111111", 
 "111111111111111100001111111111111111110000001110000001111111111111000000111111111111111111", 
 "111111111111111100000000000000111111000000001110000011100000000111000000001111111111111111", 
 "111111111111111100000000000000111110000000001110001111100000000011111000001111111111111111", 
 "111111111111111100000000000000111110000000001110000111100000000011111000001111111111111111", 
 "111111111111111110000000000000111110000000001110000000000000000011111000001111111111111111", 
 "111111111111111111100000000000111110000000001110000000000000000011111000001111111111111111", 
 "111111111111111111100000000000111110000000001110000000000000000011111000001111111111111111", 
 "111111111111111111111111100011111000000001111111110000000011111111000000001111111111111111", 
 "111111111111111111111111100011110000000001111111100000000011111111000000001111111111111111", 
 "111111111111111111111111000011110000000001111111100000000001111111000000001111111111111111", 
 "111111111111111111111100000011110000000001111110000000000000000011111000001111111111111111", 
 "111111111111111111111100000011110000000001111110000000000000000011111000001111111111111111", 
 "111111111111111111111100000111000000000001111110000000000000000011111000001111111111111111", 
 "111111111111111111111100011111000000000111111110001111100000000011111000001111111111111111", 
 "111111111111111111111100011111000000000111111110001111100000000011110000001111111111111111", 
 "111111111111111111111100011111000000000111111110000011111111111111000000001111111111111111", 
 "111111111111111111111100011111000000000111111110000001111111111111000000001111111111111111", 
 "111111111111111111111100000000000000111111111110000001111111111111000000001111111111111111", 
 "111111111111111111111100000000000000111111111111100000000000000000000000001111111111111111", 
 "111111111111111111111100000000000000111111111111100000000000000000000000001111111111111111", 
 "111111111111111111111100000000000000111111111111110000000000000000000000001111111111111111", 
 "111111111111111111111111100000000000111111111111111100000000000000000000111111111111111111", 
 "111111111111111111111111100000000000111111111111111100000000000000000000111111111111111111", 
 "111111111111111111111111100000000001111111111111111110000000000000000001111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




seventy_four <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111110000000000000000000000001111111111111111100000000000111111111111111111111", 
 "111111111111111100000000000000000000000001111111111111111100000000000111111111111111111111", 
 "111111111111111100000000000000000000000000111111111111111000000000000111111111111111111111", 
 "111111111111111100000010000000000000000000001111111111100000000000000000111111111111111111", 
 "111111111111111100001111111111111111110000001111111111100000011111000000111111111111111111", 
 "111111111111111100001111111111111111110000001111111111100000011111000000111111111111111111", 
 "111111111111111100000000000000111110000000001111111100000011111111000000111111111111111111", 
 "111111111111111100000000000000111110000000001111111100000011111111000000111111111111111111", 
 "111111111111111110000000000000111110000000001111110000000011111111000000111111111111111111", 
 "111111111111111111100000000000111110000000001111100000001111111111000000111111111111111111", 
 "111111111111111111100000000000111110000000001111100000011111111111000000111111111111111111", 
 "111111111111111111111111000011111000000001111110000001111100011111000000111111111111111111", 
 "111111111111111111111111100011110000000001111110000001111100011111000000111111111111111111", 
 "111111111111111111111111000011110000000001111110000001111000011111000000111111111111111111", 
 "111111111111111111111100000011110000000001111110001111100000011111000000111111111111111111", 
 "111111111111111111111100000011110000000001111110001111100000011111000000111111111111111111", 
 "111111111111111111111100000111000000000001111110001111100000111111000000001111111111111111", 
 "111111111111111111111100011111000000000111111110001111111111111111111000001111111111111111", 
 "111111111111111111111100011111000000000111111110001111111111111111110000001111111111111111", 
 "111111111111111111111100011111000000000111111110000000000000011111000000001111111111111111", 
 "111111111111111111111100011111000000000111111110000000000000011111000000001111111111111111", 
 "111111111111111111111100000000000000001111111110000000000000011110000000001111111111111111", 
 "111111111111111111111100000000000000111111111111100000000000000000000000001111111111111111", 
 "111111111111111111111100000000000000111111111111100000000000000000000000001111111111111111", 
 "111111111111111111111100000000000000111111111111110000000000000000000000001111111111111111", 
 "111111111111111111111111000000000000111111111111111111111111000000000000111111111111111111", 
 "111111111111111111111111100000000000111111111111111111111111000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




seventy_five <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111000000000000000000000000011111110000000000000000000000000001111111111111111", 
 "111111111111111000000000000000000000000011111110000000000000000000000000001111111111111111", 
 "111111111111111000000000000000000000000000111110000000000000000000000000001111111111111111", 
 "111111111111111000111111111111111111000000111110000111111111111111110000001111111111111111", 
 "111111111111111000111111111111111111000000111110001111111111111111111000001111111111111111", 
 "111111111111111000000000000001111100000000111110001111100000000000000000001111111111111111", 
 "111111111111111000000000000001111100000000111110001111100000000000000000001111111111111111", 
 "111111111111111000000000000001111100000000111110001111100000000000000000001111111111111111", 
 "111111111111111110000000000001111100000000111110001111111111111110000000001111111111111111", 
 "111111111111111111000000000001111100000000111110001111111111111111000000001111111111111111", 
 "111111111111111111000000000001110000000000111110000010000000000111000000001111111111111111", 
 "111111111111111111111110000111100000000011111110000000000000000011111000001111111111111111", 
 "111111111111111111111110000111100000000011111110000000000000000011111000001111111111111111", 
 "111111111111111111111000000111100000000011111110000000000000000011111000001111111111111111", 
 "111111111111111111110000000111100000000011111110000000000000000011111000001111111111111111", 
 "111111111111111111110000001111100000000011111110000000000000000011111000001111111111111111", 
 "111111111111111111110000111100000000011111111110000111100000000011111000001111111111111111", 
 "111111111111111111110000111100000000011111111110001111100000000011111000001111111111111111", 
 "111111111111111111110000111100000000011111111110000111100000000111110000001111111111111111", 
 "111111111111111111110000111100000000011111111110000001111111111111000000001111111111111111", 
 "111111111111111111110000111100000000011111111110000001111111111111000000001111111111111111", 
 "111111111111111111110000000000000011111111111110000000000000000000000000001111111111111111", 
 "111111111111111111110000000000000011111111111111100000000000000000000000001111111111111111", 
 "111111111111111111110000000000000011111111111111100000000000000000000000001111111111111111", 
 "111111111111111111111000000000000011111111111111111000000000000000000000011111111111111111", 
 "111111111111111111111110000000000011111111111111111100000000000000000000111111111111111111", 
 "111111111111111111111110000000000011111111111111111100000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




seventy_six  <=

("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111100000000000000000000000011111111111110000000000000111111111111111111111111", 
 "111111111111111100000000000000000000000001111111111100000000000000111111111111111111111111", 
 "111111111111111100000000000000000000000000111111111100000000000000011111111111111111111111", 
 "111111111111111100000100000000000001000000011111110000000000000000000111111111111111111111", 
 "111111111111111100011111111111111111100000011111110000001111111000000111111111111111111111", 
 "111111111111111100000000000001111110000000011111000000001110000000000111111111111111111111", 
 "111111111111111100000000000000111110000000011110000001111100000000000111111111111111111111", 
 "111111111111111100000000000000111110000000011110000001111100000000000111111111111111111111", 
 "111111111111111110000000000000111110000000011110000011100000000000000111111111111111111111", 
 "111111111111111111100000000000111110000000011110000111100000000000000111111111111111111111", 
 "111111111111111111100000000000111110000000011110000111100000000000000111111111111111111111", 
 "111111111111111111111111000111110000000001111110001111111111111111000000111111111111111111", 
 "111111111111111111111111000011110000000001111110000111111111111111000000111111111111111111", 
 "111111111111111111111100000011110000000001111110000111110000000111000000001111111111111111", 
 "111111111111111111111000000011110000000001111110000111100000000011111000000111111111111111", 
 "111111111111111111111000000011110000000001111110000111100000000011111000000111111111111111", 
 "111111111111111111111000000110000000000011111110000111100000000011111000000111111111111111", 
 "111111111111111111111000011110000000001111111110000111100000000011111000000111111111111111", 
 "111111111111111111111100011110000000001111111110000111100000000011111000000111111111111111", 
 "111111111111111111111000011110000000001111111110000001111111111111000000001111111111111111", 
 "111111111111111111111000011110000000001111111110000001111111111111000000000111111111111111", 
 "111111111111111111111000000000000001011111111110000001111111111111000000000111111111111111", 
 "111111111111111111111000000000000001111111111111110000000000000000000000000111111111111111", 
 "111111111111111111111000000000000001111111111111110000000000000000000000000111111111111111", 
 "111111111111111111111100000000000001111111111111110000000000000000000000001111111111111111", 
 "111111111111111111111111000000000001111111111111111100000000000000000000111111111111111111", 
 "111111111111111111111111000000000001111111111111111100000000000000000000111111111111111111", 
 "111111111111111111111111100000000001111111111111111110000111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




seventy_seven<=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111100000000000000000000000001111111000000000000000000000000111111111111111111", 
 "111111111111111100000000000000000000000001111111000000000000000000000000011111111111111111", 
 "111111111111111100000000000000000000000001111111000000000000000000000000011111111111111111", 
 "111111111111111100000000000000000000000000011111000000000000000000000000000111111111111111", 
 "111111111111111100011111111111111111100000011111000111111111111111111100000111111111111111", 
 "111111111111111100001111111111111111100000011111000011111111111111111000000111111111111111", 
 "111111111111111100000000000000111110000000011111000000000000001111100000000111111111111111", 
 "111111111111111100000000000000111110000000011111000000000000001111100000000111111111111111", 
 "111111111111111110000000000000111110000000011111000000000000001111100000000111111111111111", 
 "111111111111111111100000000000111110000000011111110000000000001111100000000111111111111111", 
 "111111111111111111100000000000111110000000011111111000000000001111000000000111111111111111", 
 "111111111111111111111111000011110000000001111111111111110000111100000000011111111111111111", 
 "111111111111111111111111000011110000000001111111111111110001111100000000011111111111111111", 
 "111111111111111111111111000011110000000001111111111111110001111100000000011111111111111111", 
 "111111111111111111111000000011110000000001111111111110000001111100000000011111111111111111", 
 "111111111111111111111000000011110000000001111111111110000001111100000000011111111111111111", 
 "111111111111111111111000000110000000000011111111111110000001100000000000111111111111111111", 
 "111111111111111111111000011110000000001111111111111110000111100000000011111111111111111111", 
 "111111111111111111111000011110000000001111111111111110001111100000000011111111111111111111", 
 "111111111111111111111000011110000000001111111111111110001111100000000011111111111111111111", 
 "111111111111111111111000011110000000001111111111111110000111100000000011111111111111111111", 
 "111111111111111111111000000000000000001111111111111110000000000000000011111111111111111111", 
 "111111111111111111111000000000000001111111111111111110000000000000011111111111111111111111", 
 "111111111111111111111000000000000001111111111111111110000000000000011111111111111111111111", 
 "111111111111111111111100000000000001111111111111111111000000000000011111111111111111111111", 
 "111111111111111111111111000000000001111111111111111111110000000000011111111111111111111111", 
 "111111111111111111111111000000000001111111111111111111110000000000011111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




seventy_eight<=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111110000100000000000001000011111111111010000000000000100111111111111111111111", 
 "111111111111111100000000000000000000000001111111110000000000000000000111111111111111111111", 
 "111111111111111100000000000000000000000001111111110000000000000000000111111111111111111111", 
 "111111111111111100000000000000000000000000011110000000000000000000000000111111111111111111", 
 "111111111111111100011111111111111111100000011110000001111111111111000000111111111111111111", 
 "111111111111111100011111111111111111100000011110000111100000000011111000001111111111111111", 
 "111111111111111100000000000000111110000000011110000111100000000011111000000111111111111111", 
 "111111111111111100000000000000111110000000011110000111100000000011111000000111111111111111", 
 "111111111111111100000000000000111110000000011110000111110000000011111000000111111111111111", 
 "111111111111111111000000000000111110000000011110000111111100000011111000000111111111111111", 
 "111111111111111111100000000000111110000000011110000111111100000011111000000111111111111111", 
 "111111111111111111100000000001110000000000011110000001111110000111000000001111111111111111", 
 "111111111111111111111111000011110000000001111110000001111111111111000000000111111111111111", 
 "111111111111111111111111000011110000000001111110000001111111111111000000000111111111111111", 
 "111111111111111111111000000011110000000001111110000111100000011111111000000111111111111111", 
 "111111111111111111111000000011110000000001111110000111100000011111111000000111111111111111", 
 "111111111111111111111000000111000000000001111110000111100000000111111000000111111111111111", 
 "111111111111111111111000011110000000001111111110000111100000000011111000000111111111111111", 
 "111111111111111111111000011110000000001111111110000111100000000011111000000111111111111111", 
 "111111111111111111111000011110000000001111111110000011110000000111000000001111111111111111", 
 "111111111111111111111000011110000000001111111110000001111111111111000000000111111111111111", 
 "111111111111111111111000000000000000001111111110000001111111111111000000000111111111111111", 
 "111111111111111111111000000000000001111111111111000000000000000000000000000111111111111111", 
 "111111111111111111111000000000000001111111111111110000000000000000000000000111111111111111", 
 "111111111111111111111000000000000001111111111111110000000000000000000000001111111111111111", 
 "111111111111111111111111000000000001111111111111111100000000000000000000111111111111111111", 
 "111111111111111111111111000000000001111111111111111100000000000000000000111111111111111111", 
 "111111111111111111111111100000000001111111111111111110000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




seventy_nine <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111100000000000000000000000001111111111000000000000000000011111111111111111111", 
 "111111111111111100000000000000000000000001111111110000000000000000000011111111111111111111", 
 "111111111111111100000000000000000000000001111111110000000000000000000011111111111111111111", 
 "111111111111111100000100000000000001000000011111000000000000000000000000011111111111111111", 
 "111111111111111100011111111111111111100000011111000000111111111111100000011111111111111111", 
 "111111111111111100000000000000111110000000011111000001110000000011100000000111111111111111", 
 "111111111111111100000000000000111110000000011111000111110000000001111100000111111111111111", 
 "111111111111111100000000000000111110000000011111000111110000000001111100000111111111111111", 
 "111111111111111111000000000000111110000000011111000111110000000001111100000111111111111111", 
 "111111111111111111100000000000111110000000011111000111110000000001111100000111111111111111", 
 "111111111111111111100000000000111110000000011111000111110000000001111100000111111111111111", 
 "111111111111111111111111000111110000000001111111000001111111111111111100000111111111111111", 
 "111111111111111111111111000011110000000001111111000000111111111111111100000111111111111111", 
 "111111111111111111111111000011110000000001111111000000111111111111111100000111111111111111", 
 "111111111111111111111000000011110000000001111111110000000000000001111100000111111111111111", 
 "111111111111111111111000000111110000000001111111111000000000000001111000000111111111111111", 
 "111111111111111111111000000110000000000011111111111000000000000011100000000111111111111111", 
 "111111111111111111111000011110000000001111111111111110000000001111100000000111111111111111", 
 "111111111111111111111000011110000000001111111111111110000000001111000000000111111111111111", 
 "111111111111111111111000011110000000001111111111111110000111111100000000000111111111111111", 
 "111111111111111111111000011110000000001111111111111110000111111100000000000111111111111111", 
 "111111111111111111111000000000000001111111111111111110000111111100000000000111111111111111", 
 "111111111111111111111000000000000001111111111111111110000000000000000000011111111111111111", 
 "111111111111111111111000000000000001111111111111111110000000000000000000011111111111111111", 
 "111111111111111111111100000000000001111111111111111111000000000000000000111111111111111111", 
 "111111111111111111111111000000000001111111111111111111110000000000000011111111111111111111", 
 "111111111111111111111111000000000001111111111111111111110000000000000011111111111111111111", 
 "111111111111111111111111100000000011111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");





eighty       <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111100000000000000000011111111111111001000000000000000111111111111111111111", 
 "111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111", 
 "111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111", 
 "111111111111111100000000000000000000000001111111000000000000000000000000111111111111111111", 
 "111111111111111100000011111111111110000001111111000001111111111111000000011111111111111111", 
 "111111111111111100011111000000001111100000011111000001111000000111100000001111111111111111", 
 "111111111111111100011111000000000111100000011111000111110000000011111000000111111111111111", 
 "111111111111111100011111000000000111100000011111000111110000000011111000000111111111111111", 
 "111111111111111100011111100000000111100000011111000111110000000011111000000111111111111111", 
 "111111111111111100011111111000000111100000011111000111110000001111111000000111111111111111", 
 "111111111111111100011111111000000111100000011111000111110000001111111000000111111111111111", 
 "111111111111111100000011111111111110000000011111000111110001100011111000000111111111111111", 
 "111111111111111100000011111111111110000000011111000111110001100011111000000111111111111111", 
 "111111111111111100000011111111111110000000011111000111110000100011111000000111111111111111", 
 "111111111111111100011111000000111111100000011111000111111100000011111000000111111111111111", 
 "111111111111111100011111000000111111100000011111000111111100000011111000000111111111111111", 
 "111111111111111100011111000000001111100000011111000111110000000011111000000111111111111111", 
 "111111111111111100011111000000000111100000011111000111110000000011111000000111111111111111", 
 "111111111111111100011111000000000111100000011111000111110000000011111000000111111111111111", 
 "111111111111111100000111111111111110000000011111000001111111111111100000000111111111111111", 
 "111111111111111100000011111111111110000000011111000001111111111111000000000111111111111111", 
 "111111111111111100000011111111111100000000011111000001111111111111000000000111111111111111", 
 "111111111111111111000000000000000000000000011111110000000000000000000000000111111111111111", 
 "111111111111111111000000000000000000000000011111110000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000011111111000000000000000000000000111111111111111", 
 "111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111", 
 "111111111111111111111000000000000000000001111111111110000000000000000000011111111111111111", 
 "111111111111111111111100000000000000000011111111111111000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




eighty_one   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111110000000000011111111111111111111111", 
 "111111111111111111100000000000000000000111111111111111110000000000011111111111111111111111", 
 "111111111111111111100000000000000000000111111111111110000000000000000111111111111111111111", 
 "111111111111111110000000000000000000000001111111111110000001111000000111111111111111111111", 
 "111111111111111110000001111111111111000000111111111110000001111100000111111111111111111111", 
 "111111111111111110000011100000000111000000001111111110000001111100000111111111111111111111", 
 "111111111111111110001111100000000011110000001111111110001111111100000111111111111111111111", 
 "111111111111111110001111100000000011110000001111111110001011111100000111111111111111111111", 
 "111111111111111110001111110000000011110000001111111110000001111100000111111111111111111111", 
 "111111111111111110001111111000000011110000001111111110000001111100000111111111111111111111", 
 "111111111111111110001111111100000011110000001111111110000001111100000111111111111111111111", 
 "111111111111111110000011111111111111000000001111111111110001111100000111111111111111111111", 
 "111111111111111110000001111111111111000000001111111111110001111100000111111111111111111111", 
 "111111111111111110000001111111111111000000001111111111110001111100000111111111111111111111", 
 "111111111111111110001111100000011111110000001111111111110001111100000111111111111111111111", 
 "111111111111111110001111100000011111110000001111111111100001111100000111111111111111111111", 
 "111111111111111110001111100000000111110000001111110000000001111100000000111111111111111111", 
 "111111111111111110001111100000000011110000001111110000000001111100000000111111111111111111", 
 "111111111111111110001111100000000011110000001111110000000001111100000000011111111111111111", 
 "111111111111111110000011100000000111000000001111110001111111111111111000000111111111111111", 
 "111111111111111110000001111111111111000000001111110000111111111111111000000111111111111111", 
 "111111111111111110000001111111111111000000001111110000000000000000000000000111111111111111", 
 "111111111111111110000000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000001111111000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000000111111111110000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000000111111111110000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000001111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");





eighty_two   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111110000000000000000000111111111111000000000000000000011111111111111111111", 
 "111111111111111111100000000000000000000111111111111000000000000000000011111111111111111111", 
 "111111111111111110000000000000000000000001111111000000000000000000000000111111111111111111", 
 "111111111111111110000001111111111110000000111111000000111111111111100000011111111111111111", 
 "111111111111111110000011100000000111000000001111000000111111111111100000011111111111111111", 
 "111111111111111110001111100000000011110000001111000001110000000011100000000111111111111111", 
 "111111111111111110001111100000000011110000001111000111110000000001111000000111111111111111", 
 "111111111111111110001111110000000011110000001111000111110000000001111000000111111111111111", 
 "111111111111111110001111111000000011110000001111000111110000001111111000000111111111111111", 
 "111111111111111110001111111100000011110000001111000111110000001111111000000111111111111111", 
 "111111111111111110001111111100000111110000001111000011100000001111111000000111111111111111", 
 "111111111111111110000001111111111111000000001111000000000001111111100000000111111111111111", 
 "111111111111111110000001111111111111000000001111000000000000111111100000000111111111111111", 
 "111111111111111110000011100000111111000000001111000000000001111100000000000111111111111111", 
 "111111111111111110001111100000011111110000001111111000000111111100000000000111111111111111", 
 "111111111111111110001111100000011111110000001111110000000111111100000000000111111111111111", 
 "111111111111111110001111100000000111110000001111000000111111100000000000011111111111111111", 
 "111111111111111110001111100000000011110000001111000000111111100000000000011111111111111111", 
 "111111111111111110001111100000000011110000001111000000111111100000000000011111111111111111", 
 "111111111111111110000001111111111111000000001111000111111111111111111100000111111111111111", 
 "111111111111111110000001111111111111000000001111000111111111111111111000000111111111111111", 
 "111111111111111110000000000000000000000000001111000001000000000000010000000111111111111111", 
 "111111111111111111100000000000000000000000001111000000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000001111000000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000001111100000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000000111111111000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000000111111111000000000000000000000000111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");





eighty_three <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111100000000000000000011111111111110000000000000000000111111111111111111111", 
 "111111111111111111000000000000000000001111111111110000000000000000000111111111111111111111", 
 "111111111111111111000000000000000000001111111111100000000000000000000111111111111111111111", 
 "111111111111111100000000000000000000000001111110000000000000000000000000111111111111111111", 
 "111111111111111100000011111111111110000001111110000001111111111111000000111111111111111111", 
 "111111111111111100011111000000000111100000011110000011110000000111000000001111111111111111", 
 "111111111111111100011111000000000111100000011110001111100000000011110000001111111111111111", 
 "111111111111111100011111000000000111100000011110001111100000000011110000001111111111111111", 
 "111111111111111100011111110000000111100000011110000000000000000011110000001111111111111111", 
 "111111111111111100011111111000000111100000011110000000000000000011110000001111111111111111", 
 "111111111111111100011111111000000111100000011110000000000000000011110000001111111111111111", 
 "111111111111111100000011111111111110000000011111110000000011111111000000001111111111111111", 
 "111111111111111100000011111111111110000000011111110000000001111111000000001111111111111111", 
 "111111111111111100000011111111111110000000011111100000000001111111000000001111111111111111", 
 "111111111111111100011111000000111111100000011110000000000000000011110000001111111111111111", 
 "111111111111111100011111000000111111100000011110000000000000000011110000001111111111111111", 
 "111111111111111100011111000000001111100000011110000000000000000011110000001111111111111111", 
 "111111111111111100011111000000000111100000011110001111100000000011110000001111111111111111", 
 "111111111111111100011111000000000111100000011110001111100000000011110000001111111111111111", 
 "111111111111111100000111111111111110000000011110000011111111111111000000001111111111111111", 
 "111111111111111100000011111111111110000000011110000001111111111111000000001111111111111111", 
 "111111111111111100000011111111111110000000011110000001111111111111000000001111111111111111", 
 "111111111111111111000000000000000000000000011111100000000000000000000000001111111111111111", 
 "111111111111111111000000000000000000000000011111110000000000000000000000001111111111111111", 
 "111111111111111111100000000000000000000000011111110000000000000000000000001111111111111111", 
 "111111111111111111111000000000000000000001111111111100000000000000000000111111111111111111", 
 "111111111111111111111000000000000000000001111111111100000000000000000000111111111111111111", 
 "111111111111111111111100000000000000000011111111111110000000000000000001111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");





eighty_four  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111100000000000000000001111111111111111111100000000000111111111111111111111", 
 "111111111111111111000000000000000000001111111111111111111100000000000111111111111111111111", 
 "111111111111111111000000000000000000001111111111111111111000000000000111111111111111111111", 
 "111111111111111100000000000000000000000001111111111111100000000000000000111111111111111111", 
 "111111111111111100000011111111111110000001111111111111100000011111000000111111111111111111", 
 "111111111111111100011111000000000111100000011111111111100000011111000000111111111111111111", 
 "111111111111111100011111000000000111100000011111111100000001111111000000111111111111111111", 
 "111111111111111100011111000000000111100000011111111100000011111111000000111111111111111111", 
 "111111111111111100011111100000000111100000011111110000000011111111000000111111111111111111", 
 "111111111111111100011111111000000111100000011111110000001111111111000000111111111111111111", 
 "111111111111111100011111111000001111100000011111100000001111111111000000111111111111111111", 
 "111111111111111100000111111111111110000000011110000001111100011111000000111111111111111111", 
 "111111111111111100000011111111111110000000011110000001111100011111000000111111111111111111", 
 "111111111111111100000011111111111110000000011110000001111100011111000000111111111111111111", 
 "111111111111111100011111000000111111100000011110001111100000011111000000111111111111111111", 
 "111111111111111100011111000000111111100000011110001111100000011111000000111111111111111111", 
 "111111111111111100011111000000001111100000011110001111110000111111000000001111111111111111", 
 "111111111111111100011111000000000111100000011110001111111111111111110000001111111111111111", 
 "111111111111111100011111000000000111100000011110001111111111111111110000001111111111111111", 
 "111111111111111100000111111111111110000000011110000000000000011111000000001111111111111111", 
 "111111111111111100000011111111111110000000011110000000000000011111000000001111111111111111", 
 "111111111111111100000011111111111100000000011110000000000000011111000000001111111111111111", 
 "111111111111111111000000000000000000000000011111100000000000000000000000001111111111111111", 
 "111111111111111111000000000000000000000000011111110000000000000000000000001111111111111111", 
 "111111111111111111100000000000000000000000011111110000000000000000000000001111111111111111", 
 "111111111111111111111000000000000000000001111111111111111111000000000000111111111111111111", 
 "111111111111111111111000000000000000000001111111111111111111000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");





eighty_five  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111000000000000000000001111111110000000000000000000000000001111111111111111", 
 "111111111111111111000000000000000000001111111110000000000000000000000000001111111111111111", 
 "111111111111111100000000000000000000000011111110000000000000000000000000001111111111111111", 
 "111111111111111100000011111111111100000001111110000111111111111111110000001111111111111111", 
 "111111111111111100000111000000001110000000011110001111111111111111110000001111111111111111", 
 "111111111111111100011111000000000111100000011110001111100000000000000000001111111111111111", 
 "111111111111111100011111000000000111100000011110001111100000000000000000001111111111111111", 
 "111111111111111100011111000000000111100000011110001111100000000000000000001111111111111111", 
 "111111111111111100011111110000000111100000011110001111111111111111000000001111111111111111", 
 "111111111111111100011111111000000111100000011110001111111111111111000000001111111111111111", 
 "111111111111111100000111111000001110000000011110000010000000000111000000001111111111111111", 
 "111111111111111100000011111111111110000000011110000000000000000011110000001111111111111111", 
 "111111111111111100000011111111111110000000011110000000000000000011110000001111111111111111", 
 "111111111111111100000111000001111110000000011110000000000000000011110000001111111111111111", 
 "111111111111111100011111000000111111100000011110000000000000000011110000001111111111111111", 
 "111111111111111100011111000000111111100000011110000000000000000011110000001111111111111111", 
 "111111111111111100011111000000001111100000011110000111100000000011110000001111111111111111", 
 "111111111111111100011111000000000111100000011110001111100000000011110000001111111111111111", 
 "111111111111111100001111000000001111100000011110000111100000000111110000001111111111111111", 
 "111111111111111100000011111111111110000000011110000001111111111111000000001111111111111111", 
 "111111111111111100000011111111111110000000011110000001111111111111000000001111111111111111", 
 "111111111111111100000000000000000000000000011110000000000000000000000000001111111111111111", 
 "111111111111111111000000000000000000000000011111100000000000000000000000001111111111111111", 
 "111111111111111111000000000000000000000000011111110000000000000000000000001111111111111111", 
 "111111111111111111100000000000000000000000111111111000000000000000000000011111111111111111", 
 "111111111111111111111000000000000000000001111111111100000000000000000000111111111111111111", 
 "111111111111111111111000000000000000000001111111111100000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");





eighty_six   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111110000000000000000001111111111111110000000000000111111111111111111111111", 
 "111111111111111111100000000000000000000111111111111110000000000000111111111111111111111111", 
 "111111111111111111100000000000000000000111111111111100000000000000111111111111111111111111", 
 "111111111111111110000000000000000000000000111111110000000000000000000111111111111111111111", 
 "111111111111111110000001111111111111000000111111110000001111111000000111111111111111111111", 
 "111111111111111110001111100000000011110000001111000000001110000000000111111111111111111111", 
 "111111111111111110001111100000000011110000001110000001111100000000000111111111111111111111", 
 "111111111111111110001111100000000011110000001110000001111100000000000111111111111111111111", 
 "111111111111111110001111110000000011110000001110000011110000000000000111111111111111111111", 
 "111111111111111110001111111100000011110000001110000111100000000000000111111111111111111111", 
 "111111111111111110001111111100000011110000001110000111110000000000000111111111111111111111", 
 "111111111111111110000001111111111111000000001110001111111111111111000000111111111111111111", 
 "111111111111111110000001111111111111000000001110000111111111111111000000111111111111111111", 
 "111111111111111110000001110000111111000000001110000111110000000111000000001111111111111111", 
 "111111111111111110001111100000011111110000001110000111110000000011111000001111111111111111", 
 "111111111111111110001111100000011111110000001110000111100000000011111000000111111111111111", 
 "111111111111111110001111100000000111110000001110000111100000000011111000000111111111111111", 
 "111111111111111110001111100000000011110000001110000111100000000011111000000111111111111111", 
 "111111111111111110001111100000000011110000001110000111100000000011111000000111111111111111", 
 "111111111111111110000011111111111111000000001110000001111111111111000000001111111111111111", 
 "111111111111111110000001111111111111000000001110000001111111111111000000000111111111111111", 
 "111111111111111110000001111111111110000000001110000001111111111111000000000111111111111111", 
 "111111111111111111100000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000001111110000000000000000000000001111111111111111", 
 "111111111111111111110000000000000000000000001111110000000000000000000000001111111111111111", 
 "111111111111111111111100000000000000000000111111111100000000000000000000111111111111111111", 
 "111111111111111111111100000000000000000000111111111110000000000000000000111111111111111111", 
 "111111111111111111111110000000000001100001111111111111000111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




eighty_seven <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111100000000000000000001111111110000000000000000000000001111111111111111111", 
 "111111111111111111000000000000000000001111111110000000000000000000000000111111111111111111", 
 "111111111111111111000000000000000000001111111110000000000000000000000000111111111111111111", 
 "111111111111111100000000000000000000000001111110000000000000000000000000001111111111111111", 
 "111111111111111100000011111111111110000001111110001111111111111111110000001111111111111111", 
 "111111111111111100011111000000000111100000011110000111111111111111110000001111111111111111", 
 "111111111111111100011111000000000111100000011110000000000000011111000000001111111111111111", 
 "111111111111111100011111000000000111100000011110000000000000011111000000001111111111111111", 
 "111111111111111100011111100000000111100000011111000000000000011111000000001111111111111111", 
 "111111111111111100011111111000000111100000011111110000000000011111000000001111111111111111", 
 "111111111111111100011111111000001111100000011111110000000000011111000000001111111111111111", 
 "111111111111111100000111111111111110000000011111111111100001111000000000111111111111111111", 
 "111111111111111100000011111111111110000000011111111111100001111000000000111111111111111111", 
 "111111111111111100000011111111111110000000011111111111100001111000000000111111111111111111", 
 "111111111111111100011111000000111111100000011111111100000001111000000000111111111111111111", 
 "111111111111111100011111000000111111100000011111111100000001111000000000111111111111111111", 
 "111111111111111100011111000000001111100000011111111100000011000000000001111111111111111111", 
 "111111111111111100011111000000000111100000011111111100001111000000000111111111111111111111", 
 "111111111111111100011111000000000111100000011111111100001111000000000111111111111111111111", 
 "111111111111111100000111111111111110000000011111111100001111000000000111111111111111111111", 
 "111111111111111100000011111111111110000000011111111100001111000000000111111111111111111111", 
 "111111111111111100000011111111111100000000011111111100000000000000000111111111111111111111", 
 "111111111111111111000000000000000000000000011111111100000000000000111111111111111111111111", 
 "111111111111111111000000000000000000000000011111111100000000000000111111111111111111111111", 
 "111111111111111111100000000000000000000000011111111110000000000000111111111111111111111111", 
 "111111111111111111111000000000000000000001111111111111100000000000111111111111111111111111", 
 "111111111111111111111000000000000000000001111111111111100000000000111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");





eighty_eight <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111110010000000000000101111111111111000000000000000100111111111111111111111", 
 "111111111111111111100000000000000000000111111111110000000000000000000111111111111111111111", 
 "111111111111111111100000000000000000000111111111110000000000000000000111111111111111111111", 
 "111111111111111110000000000000000000000001111110000000000000000000000000111111111111111111", 
 "111111111111111110000001111111111110000000111110000001111111111111000000111111111111111111", 
 "111111111111111110001111100000000111110000001110000111110000000011110000001111111111111111", 
 "111111111111111110001111100000000011110000001110000111100000000011111000000111111111111111", 
 "111111111111111110001111100000000011110000001110000111110000000011111000000111111111111111", 
 "111111111111111110001111110000000011110000001110000111110000000011111000000111111111111111", 
 "111111111111111110001111111000000011110000001110000111111100000011111000000111111111111111", 
 "111111111111111110001111111100000011110000001110000111111100000011111000001111111111111111", 
 "111111111111111110000011111100000111000000001110000001111110000111000000001111111111111111", 
 "111111111111111110000001111111111111000000001110000001111111111111000000001111111111111111", 
 "111111111111111110000001111111111111000000001110000001111111111111000000000111111111111111", 
 "111111111111111110001111100000011111110000001110000111110000011111110000000111111111111111", 
 "111111111111111110001111100000011111110000001110000111100000011111111000000111111111111111", 
 "111111111111111110001111100000000111110000001110000111100000000111111000000111111111111111", 
 "111111111111111110001111100000000011110000001110000111100000000011111000000111111111111111", 
 "111111111111111110001111100000000011110000001110000111100000000011111000000111111111111111", 
 "111111111111111110000011100000000111000000001110000011110000000111000000001111111111111111", 
 "111111111111111110000001111111111111000000001110000001111111111111000000001111111111111111", 
 "111111111111111110000001111111111111000000001110000001111111111111000000000111111111111111", 
 "111111111111111110000000000000000000000000001111000000000000000000000000000111111111111111", 
 "111111111111111111100000000000000000000000001111110000000000000000000000000111111111111111", 
 "111111111111111111110000000000000000000000001111110000000000000000000000001111111111111111", 
 "111111111111111111111100000000000000000000111111111100000000000000000000111111111111111111", 
 "111111111111111111111100000000000000000000111111111110000000000000000000111111111111111111", 
 "111111111111111111111110000000000000000001111111111110000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




eighty_nine  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111100000000000000000001111111111110000000000000000000111111111111111111111", 
 "111111111111111111000000000000000000001111111111110000000000000000000111111111111111111111", 
 "111111111111111111000000000000000000001111111111100000000000000000000111111111111111111111", 
 "111111111111111100000000000000000000000001111110000000000000000000000000111111111111111111", 
 "111111111111111100000011100000011110000000111110000001111111111111000000111111111111111111", 
 "111111111111111100011111000000000111100000011110000011110000000111000000001111111111111111", 
 "111111111111111100011111000000000111100000011110001111100000000011110000001111111111111111", 
 "111111111111111100011111000000000111100000011110001111100000000011110000001111111111111111", 
 "111111111111111100011111110000000111100000011110001111100000000011110000001111111111111111", 
 "111111111111111100011111111000000111100000011110001111100000000011110000001111111111111111", 
 "111111111111111100011111111000000111100000011110001111100000000011111000001111111111111111", 
 "111111111111111100000011111111111110000000011110000001111111111111111000001111111111111111", 
 "111111111111111100000011111111111110000000011110000001111111111111110000001111111111111111", 
 "111111111111111100000011111111111110000000011110000001111111111111110000001111111111111111", 
 "111111111111111100011111000000111111100000011111110000000000000011110000001111111111111111", 
 "111111111111111100011111000000111111100000011111110000000000000011110000001111111111111111", 
 "111111111111111100011111000000001111100000011111110000000000000111000000001111111111111111", 
 "111111111111111100011111000000000111100000011111111100000000011111000000001111111111111111", 
 "111111111111111100011111000000000111100000011111111100000000011111000000001111111111111111", 
 "111111111111111100000111111111111110000000011111111100001111111000000000001111111111111111", 
 "111111111111111100000011111111111110000000011111111100001111111000000000001111111111111111", 
 "111111111111111100000011111111111100000000011111111100001111111000000000001111111111111111", 
 "111111111111111111000000000000000000000000011111111100000000000000000000111111111111111111", 
 "111111111111111111000000000000000000000000011111111100000000000000000000111111111111111111", 
 "111111111111111111100000000000000000000000011111111110000000000000000001111111111111111111", 
 "111111111111111111111000000000000000000001111111111111100000000000000111111111111111111111", 
 "111111111111111111111000000000000000000001111111111111100000000000000111111111111111111111", 
 "111111111111111111111110000000000011000111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




ninety       <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111100000000000000000011111111111111100000000000000000011111111111111111111", 
 "111111111111111111000000000000000000001111111111111000000000000000000011111111111111111111", 
 "111111111111111111000000000000000000001111111111110000000000000000000001111111111111111111", 
 "111111111111111100000000000000000000000011111111000000000000000000000000011111111111111111", 
 "111111111111111100000111111111111100000011111111000000111111111111100000011111111111111111", 
 "111111111111111100000111100000011110000000111111000000111000000011100000000111111111111111", 
 "111111111111111100011111000000001111100000011111000011111000000001111100000111111111111111", 
 "111111111111111100011111000000001111100000011111000011110000000001111100000111111111111111", 
 "111111111111111100011111000000001111100000011111000011110000000011111100000111111111111111", 
 "111111111111111100011111000000001111100000011111000011110000001111111100000111111111111111", 
 "111111111111111100011111000000001111100000011111000011111000001111111100000111111111111111", 
 "111111111111111100000111111111111111100000011111000111111000110001111100000111111111111111", 
 "111111111111111100000111111111111111100000011111000011110000110001111100000111111111111111", 
 "111111111111111100000011111111111111100000011111000011111000100001111100000111111111111111", 
 "111111111111111111000000000000001111100000011111000011111110000001111100000111111111111111", 
 "111111111111111111000000000000001111100000011111000011111110000001111100000111111111111111", 
 "111111111111111111100000000000001110000000011111000011111000000001111100000111111111111111", 
 "111111111111111111111000000001111100000000011111000011111000000001111100000111111111111111", 
 "111111111111111111111000000001111100000000011111000011110000000001111100000111111111111111", 
 "111111111111111111111000111111110000000000011111000000111111111111100000000111111111111111", 
 "111111111111111111111000111111110000000000011111000000111111111111100000000111111111111111", 
 "111111111111111111111000011111100000000000011111000000111111111111100000000111111111111111", 
 "111111111111111111111000000000000000000001111111111000000000000000000000000111111111111111", 
 "111111111111111111111000000000000000000011111111111000000000000000000000000111111111111111", 
 "111111111111111111111000000000000000000011111111111000000000000000000000000111111111111111", 
 "111111111111111111111111000000000000001111111111111111000000000000000000011111111111111111", 
 "111111111111111111111111000000000000011111111111111111000000000000000000011111111111111111", 
 "111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




ninety_one   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111000000000000000000001111111111111111100000000000111111111111111111111111", 
 "111111111111111111000000000000000000001111111111111111100000000000011111111111111111111111", 
 "111111111111111100000000000000000000000011111111111110000000000000000111111111111111111111", 
 "111111111111111100000111111111111100000011111111111100000001111000000111111111111111111111", 
 "111111111111111100000111111111111100000001111111111100000001111000000111111111111111111111", 
 "111111111111111100000111000000001110000000011111111100000011111000000111111111111111111111", 
 "111111111111111100011111000000001111100000011111111100001111111000000111111111111111111111", 
 "111111111111111100011111000000001111100000011111111100000011111000000111111111111111111111", 
 "111111111111111100011111000000001111100000011111111100000001111000000111111111111111111111", 
 "111111111111111100011111000000001111100000011111111100000001111000000111111111111111111111", 
 "111111111111111100000111000000001111100000011111111110000001111000000111111111111111111111", 
 "111111111111111100000111111111111111100000011111111111100001111000000111111111111111111111", 
 "111111111111111100000111111111111111100000011111111111100001111000000111111111111111111111", 
 "111111111111111100000000000000001111100000011111111111100001111000000111111111111111111111", 
 "111111111111111111000000000000001111100000011111111111100001111000000111111111111111111111", 
 "111111111111111111000000000000001111100000011111111111100001111000000111111111111111111111", 
 "111111111111111111110000000000111100000000011111110000000001111000000000111111111111111111", 
 "111111111111111111111000000001111100000000011111110000000001111000000000111111111111111111", 
 "111111111111111111111000000001111100000000011111110000000011111000000000111111111111111111", 
 "111111111111111111111000111111110000000000011111110001111111111111111000000111111111111111", 
 "111111111111111111111000111111110000000000011111110001111111111111111000000111111111111111", 
 "111111111111111111111000000000000000000000011111110000000000000000000000000111111111111111", 
 "111111111111111111111000000000000000000001111111110000000000000000000000000111111111111111", 
 "111111111111111111111000000000000000000011111111110000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000111111111111000000000000000000000000111111111111111", 
 "111111111111111111111111000000000000001111111111111100000000000000000000000111111111111111", 
 "111111111111111111111111111111111111111111111111111100000000000000000000000111111111111111", 
 "111111111111111111111111111111111111111111111111111111000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




ninety_two   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111", 
 "111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111", 
 "111111111111111100000000000000000000000011111111000000000000000000000000111111111111111111", 
 "111111111111111100000011111111111100000011111110000001111111111111000000111111111111111111", 
 "111111111111111100000111111111111100000011111110000001111111111111000000111111111111111111", 
 "111111111111111100000111000000001110000000011110000001110000000011100000000111111111111111", 
 "111111111111111100011111000000001111100000011110000111110000000011111000000111111111111111", 
 "111111111111111100011111000000001111100000011110000111110000000011111000000111111111111111", 
 "111111111111111100011111000000001111100000011110000111110000001111111000000111111111111111", 
 "111111111111111100011111000000001111100000011110000111110000001111111000000111111111111111", 
 "111111111111111100011111000000001111100000011110000011100000011111110000000111111111111111", 
 "111111111111111100000111111111111111100000011110000000000001111111000000000111111111111111", 
 "111111111111111100000111111111111111100000011110000000000001111111000000000111111111111111", 
 "111111111111111100000000000000001111100000011111000000000001111100000000000111111111111111", 
 "111111111111111111000000000000001111100000011111110000001111111000000000000111111111111111", 
 "111111111111111111000000000000001111100000011111110000001111111000000000000111111111111111", 
 "111111111111111111110000000000111100000000011111000001111111100000000000011111111111111111", 
 "111111111111111111111000000001111100000000011110000001111111100000000000111111111111111111", 
 "111111111111111111111000000001111100000000011110000001111111100000000000011111111111111111", 
 "111111111111111111111000111111110000000000011111000111111111111111111000000111111111111111", 
 "111111111111111111111000111111110000000000011110000111111111111111111000000111111111111111", 
 "111111111111111111111000000000000000000000011110000001000000000000100000000111111111111111", 
 "111111111111111111111000000000000000000011111110000000000000000000000000000111111111111111", 
 "111111111111111111111000000000000000000011111110000000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000011111111000000000000000000000000000111111111111111", 
 "111111111111111111111111000000000000001111111111110000000000000000000000000111111111111111", 
 "111111111111111111111111111111111111111111111111110000000000000000000000000111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




ninety_three <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111110000000000000000001111111111111100000000000000000011111111111111111111", 
 "111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111", 
 "111111111111111111100000000000000000000111111111111000000000000000000001111111111111111111", 
 "111111111111111110000000000000000000000001111111100000100000000000000000011111111111111111", 
 "111111111111111110000011111111111110000001111111000000111111111111100000011111111111111111", 
 "111111111111111110000011100000000111000000001111000000111000000001100000000111111111111111", 
 "111111111111111110001111100000000111110000001111000011111000000001111100000011111111111111", 
 "111111111111111110001111100000000111110000001111000011111000000001111100000011111111111111", 
 "111111111111111110001111100000000111110000001111000000000000000001111100000011111111111111", 
 "111111111111111110001111100000000111110000001111000000000000000001111100000011111111111111", 
 "111111111111111110001111100000000111110000001111000000000000000001111100000011111111111111", 
 "111111111111111110000011111111111111110000001111111000000000111111100000000011111111111111", 
 "111111111111111110000011111111111111110000001111111000000000111111100000000011111111111111", 
 "111111111111111110000001111111111111110000001111111000000000111111100000000011111111111111", 
 "111111111111111111100000000000000111110000001111000000000000000001111100000011111111111111", 
 "111111111111111111100000000000000111110000001111000000000000000001111100000011111111111111", 
 "111111111111111111110000000000000111000000001111000000000000000001111100000011111111111111", 
 "111111111111111111111100000000111110000000001111000011111000000001111100000011111111111111", 
 "111111111111111111111100000000111110000000001111000011111000000001111100000011111111111111", 
 "111111111111111111111100001111111000000000001111100000111111111111110000000011111111111111", 
 "111111111111111111111100011111111000000000001111000000111111111111100000000011111111111111", 
 "111111111111111111111100011111111000000000001111000000111111111111100000000011111111111111", 
 "111111111111111111111100000000000000000000111111111000000000000000000000000011111111111111", 
 "111111111111111111111100000000000000000001111111111000000000000000000000000011111111111111", 
 "111111111111111111111100000000000000000001111111111100000000000000000000000111111111111111", 
 "111111111111111111111111100000000000000111111111111111000000000000000000011111111111111111", 
 "111111111111111111111111100000000000001111111111111111000000000000000000011111111111111111", 
 "111111111111111111111111111111111111111111111111111111100000000000000000011111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




ninety_four  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111100000000000000000011111111111111111111110000000000111111111111111111111", 
 "111111111111111111000000000000000000001111111111111111111100000000000011111111111111111111", 
 "111111111111111111000000000000000000001111111111111111111100000000000011111111111111111111", 
 "111111111111111100000000000000000000000011111111111111110000000000000000111111111111111111", 
 "111111111111111100000111111111111100000011111111111111110000001111000000111111111111111111", 
 "111111111111111100000111111111111100000001111111111111100000011111000000111111111111111111", 
 "111111111111111100011111000000001111100000011111111110000001111111000000111111111111111111", 
 "111111111111111100011111000000001111100000011111111110000001111111000000111111111111111111", 
 "111111111111111100011111000000001111100000011111110000000011111111000000111111111111111111", 
 "111111111111111100011111000000001111100000011111110000001111111111000000111111111111111111", 
 "111111111111111100011111000000001111100000011111110000001111111111000000111111111111111111", 
 "111111111111111100000111111111111111100000011111000001111100011111000000111111111111111111", 
 "111111111111111100000111111111111111100000011110000001111100011111000000111111111111111111", 
 "111111111111111100000011111111111111100000011110000001111100001111000000111111111111111111", 
 "111111111111111111000000000000001111100000011110000111110000001111000000111111111111111111", 
 "111111111111111111000000000000001111100000011110000111110000001111000000111111111111111111", 
 "111111111111111111100000000000001110000000011110000111110000011111100000000111111111111111", 
 "111111111111111111111000000001111100000000011110000111111111111111111000000111111111111111", 
 "111111111111111111111000000001111100000000011110000111111111111111111000000111111111111111", 
 "111111111111111111111000011111110000000000011111000000000000011111100000000111111111111111", 
 "111111111111111111111000111111110000000000011110000000000000001111000000000111111111111111", 
 "111111111111111111111000011111100000000000011110000000000000001111000000000111111111111111", 
 "111111111111111111111000000000000000000001111111100000000000000000000000000111111111111111", 
 "111111111111111111111000000000000000000011111111110000000000000000000000000111111111111111", 
 "111111111111111111111000000000000000000011111111110000000000000000000000001111111111111111", 
 "111111111111111111111111000000000000001111111111111111111111100000000000011111111111111111", 
 "111111111111111111111111000000000000011111111111111111111111100000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




ninety_five  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111000000000000000000001111111110000000000000000000000000000111111111111111", 
 "111111111111111111000000000000000000001111111110000000000000000000000000000111111111111111", 
 "111111111111111100000000000000000000000011111110000000000000000000000000000111111111111111", 
 "111111111111111100000011111111111100000011111110000111111111111111111000000111111111111111", 
 "111111111111111100000111111111111100000011111110000111111111111111111000000111111111111111", 
 "111111111111111100000111000000001110000000011110000111110000000000000000000111111111111111", 
 "111111111111111100011111000000001111100000011110000111110000000000000000000111111111111111", 
 "111111111111111100011111000000001111100000011110000111110000000000000000000111111111111111", 
 "111111111111111100011111000000001111100000011110000111111111111111000000000111111111111111", 
 "111111111111111100011111000000001111100000011110000111111111111111000000000111111111111111", 
 "111111111111111100000111000000001111100000011111000001000000000111100000000111111111111111", 
 "111111111111111100000111111111111111100000011110000000000000000011111000000111111111111111", 
 "111111111111111100000111111111111111100000011110000000000000000011111000000111111111111111", 
 "111111111111111100000000000000001111100000011110000000000000000011111000000111111111111111", 
 "111111111111111111000000000000001111100000011110000000000000000011111000000111111111111111", 
 "111111111111111111000000000000001111100000011110000000000000000011111000000111111111111111", 
 "111111111111111111110000000000111100000000011110000111100000000011111000000111111111111111", 
 "111111111111111111111000000001111100000000011110000111110000000011111000000111111111111111", 
 "111111111111111111111000000001111100000000011110000011110000000011110000000111111111111111", 
 "111111111111111111111000111111110000000000011110000001111111111111000000000111111111111111", 
 "111111111111111111111000111111110000000000011110000001111111111111000000000111111111111111", 
 "111111111111111111111000000000000000000000011111000000000000000000000000000111111111111111", 
 "111111111111111111111000000000000000000001111111110000000000000000000000000111111111111111", 
 "111111111111111111111000000000000000000011111111110000000000000000000000000111111111111111", 
 "111111111111111111111100000000000000000111111111111000000000000000000000001111111111111111", 
 "111111111111111111111111000000000000001111111111111110000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111110000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




ninety_six   <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111100000000000000000011111111111111110000000000000111111111111111111111111", 
 "111111111111111111000000000000000000001111111111111100000000000000111111111111111111111111", 
 "111111111111111111000000000000000000001111111111111100000000000000111111111111111111111111", 
 "111111111111111100000000000000000000000011111111100000000000000000000111111111111111111111", 
 "111111111111111100000111111111111100000011111111100000001111111000000111111111111111111111", 
 "111111111111111100000111000000001110000000011110000000011100000000000111111111111111111111", 
 "111111111111111100011111000000001111100000011110000011111100000000000111111111111111111111", 
 "111111111111111100011111000000001111100000011110000011111100000000000111111111111111111111", 
 "111111111111111100011111000000001111100000011110000011100000000000000111111111111111111111", 
 "111111111111111100011111000000001111100000011110001111100000000000000111111111111111111111", 
 "111111111111111100011111000000001111100000011110001111100000000000000111111111111111111111", 
 "111111111111111100000111111111111111100000011110001111111111111111000000111111111111111111", 
 "111111111111111100000111111111111111100000011110001111111111111111000000111111111111111111", 
 "111111111111111100000000000000011111100000011110001111110000001111000000011111111111111111", 
 "111111111111111111000000000000001111100000011110001111100000000111110000001111111111111111", 
 "111111111111111111000000000000001111100000011110001111100000000111110000001111111111111111", 
 "111111111111111111100000000000001110000000011110001111100000000111110000001111111111111111", 
 "111111111111111111111000000001111100000000011110001111100000000111110000001111111111111111", 
 "111111111111111111111000000001111100000000011110001111100000000111110000001111111111111111", 
 "111111111111111111111000111111110000000000011110000011111111111111000000001111111111111111", 
 "111111111111111111111000111111110000000000011110000011111111111111000000001111111111111111", 
 "111111111111111111111000011111100000000000011110000011111111111110000000001111111111111111", 
 "111111111111111111111000000000000000000011111111100000000000000000000000001111111111111111", 
 "111111111111111111111000000000000000000011111111100000000000000000000000001111111111111111", 
 "111111111111111111111000000000000000000011111111110000000000000000000000001111111111111111", 
 "111111111111111111111111000000000000001111111111111100000000000000000000111111111111111111", 
 "111111111111111111111111000000000000011111111111111100000000000000000001111111111111111111", 
 "111111111111111111111111111111111111111111111111111110001111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




ninety_seven <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111100000000000000000011111111111000000000000000000000000111111111111111111", 
 "111111111111111111000000000000000000001111111110000000000000000000000000111111111111111111", 
 "111111111111111111000000000000000000001111111110000000000000000000000000011111111111111111", 
 "111111111111111100000000000000000000000011111110000001000000000000000000000111111111111111", 
 "111111111111111100000111111111111100000011111110000111111111111111111000000111111111111111", 
 "111111111111111100000111111111111100000001111110000111111111111111111000000111111111111111", 
 "111111111111111100011111000000001111100000011110000000000000001111000000000111111111111111", 
 "111111111111111100011111000000001111100000011110000000000000001111000000000111111111111111", 
 "111111111111111100011111000000001111100000011111000000000000001111000000000111111111111111", 
 "111111111111111100011111000000001111100000011111110000000000001111000000000111111111111111", 
 "111111111111111100011111000000001111100000011111110000000000011111000000000111111111111111", 
 "111111111111111100000111111111111111100000011111111111100001111100000000011111111111111111", 
 "111111111111111100000111111111111111100000011111111111110001111000000000111111111111111111", 
 "111111111111111100000011111111111111100000011111111111110001111000000000111111111111111111", 
 "111111111111111111000000000000001111100000011111111110000001111000000000111111111111111111", 
 "111111111111111111000000000000001111100000011111111110000001111000000000111111111111111111", 
 "111111111111111111100000000000001110000000011111111110000001100000000000111111111111111111", 
 "111111111111111111111000000001111100000000011111111110001111100000000011111111111111111111", 
 "111111111111111111111000000001111100000000011111111110001111100000000011111111111111111111", 
 "111111111111111111111000011111110000000000011111111110001111100000000011111111111111111111", 
 "111111111111111111111000111111110000000000011111111110001111100000000011111111111111111111", 
 "111111111111111111111000011111100000000000011111111110000000000000000111111111111111111111", 
 "111111111111111111111000000000000000000001111111111110000000000000011111111111111111111111", 
 "111111111111111111111000000000000000000011111111111110000000000000011111111111111111111111", 
 "111111111111111111111000000000000000000011111111111110000000000000011111111111111111111111", 
 "111111111111111111111111000000000000001111111111111111110000000000011111111111111111111111", 
 "111111111111111111111111000000000000011111111111111111110000000000011111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");



ninety_eight <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111100100000000000010011111111111110010000000000000001111111111111111111111", 
 "111111111111111111000000000000000000001111111111100000000000000000000111111111111111111111", 
 "111111111111111111000000000000000000001111111111100000000000000000000111111111111111111111", 
 "111111111111111100000000000000000000000011111110000000000000000000000001111111111111111111", 
 "111111111111111100000111111111111100000011111110000011111111111111000000111111111111111111", 
 "111111111111111100000111111111111100000011111110000111100000000111110000001111111111111111", 
 "111111111111111100011111000000001111100000011110001111100000000111110000001111111111111111", 
 "111111111111111100011111000000001111100000011110001111100000000111110000001111111111111111", 
 "111111111111111100011111000000001111100000011110001111110000000111110000001111111111111111", 
 "111111111111111100011111000000001111100000011110001111111000000111110000001111111111111111", 
 "111111111111111100011111000000001111100000011110001111111100000111110000001111111111111111", 
 "111111111111111100000111000000001111100000011110000011111100000111000000001111111111111111", 
 "111111111111111100000111111111111111100000011110000011111111111111000000001111111111111111", 
 "111111111111111100000111111111111111100000011110000011111111111111000000001111111111111111", 
 "111111111111111111000000000000001111100000011110000111100000011111110000001111111111111111", 
 "111111111111111111000000000000001111100000011110001111100000011111110000001111111111111111", 
 "111111111111111111100000000000001110000000011110001111100000000111110000001111111111111111", 
 "111111111111111111111000000001111100000000011110001111100000000111110000001111111111111111", 
 "111111111111111111111000000001111100000000011110001111100000000111110000001111111111111111", 
 "111111111111111111111000000001110000000000011110000011100000000111000000001111111111111111", 
 "111111111111111111111000111111110000000000011110000011111111111111000000001111111111111111", 
 "111111111111111111111000111111110000000000011110000011111111111111000000001111111111111111", 
 "111111111111111111111000000000000000000000011110000000000000000000000000001111111111111111", 
 "111111111111111111111000000000000000000011111111100000000000000000000000001111111111111111", 
 "111111111111111111111000000000000000000011111111110000000000000000000000001111111111111111", 
 "111111111111111111111111000000000000001111111111111100000000000000000000111111111111111111", 
 "111111111111111111111111000000000000001111111111111100000000000000000000111111111111111111", 
 "111111111111111111111111111111111111111111111111111100000000000000000001111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




ninety_nine  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111100000000000000000011111111111110000000000000000000111111111111111111111", 
 "111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111", 
 "111111111111111111000000000000000000001111111111110000000000000000000011111111111111111111", 
 "111111111111111100000000000000000000000011111110000001000000000000000000111111111111111111", 
 "111111111111111100000111111111111100000011111110000001111111111111000000111111111111111111", 
 "111111111111111100000111000000001110000000011110000001110000000011100000001111111111111111", 
 "111111111111111100011111000000001111100000011110000111110000000011111000000111111111111111", 
 "111111111111111100011111000000001111100000011110000111110000000011111000000111111111111111", 
 "111111111111111100011111000000001111100000011110000111110000000011111000000111111111111111", 
 "111111111111111100011111000000001111100000011110000111110000000011111000000111111111111111", 
 "111111111111111100011111000000001111100000011110000111110000000011111000000111111111111111", 
 "111111111111111100000111111111111111100000011111000001111111111111111000000111111111111111", 
 "111111111111111100000111111111111111100000011110000001111111111111111000000111111111111111", 
 "111111111111111100000011111111111111100000011111000001111111111111111000000111111111111111", 
 "111111111111111111000000000000001111100000011111110000000000000011111000000111111111111111", 
 "111111111111111111000000000000001111100000011111110000000000000011111000000111111111111111", 
 "111111111111111111100000000000001110000000011111111000000000000011000000000111111111111111", 
 "111111111111111111111000000001111100000000011111111110000000001111000000000111111111111111", 
 "111111111111111111111000000001111100000000011111111110000000011111000000000111111111111111", 
 "111111111111111111111000011111110000000000011111111110001111111100000000000111111111111111", 
 "111111111111111111111000111111110000000000011111111110001111111000000000000111111111111111", 
 "111111111111111111111000011111110000000000011111111110001111111000000000000111111111111111", 
 "111111111111111111111000000000000000000011111111111110000000000000000000111111111111111111", 
 "111111111111111111111000000000000000000011111111111110000000000000000000111111111111111111", 
 "111111111111111111111000000000000000000011111111111110000000000000000000111111111111111111", 
 "111111111111111111111111000000000000001111111111111111110000000000000011111111111111111111", 
 "111111111111111111111111000000000000011111111111111111110000000000000111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");




one_hundred  <=
("111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111110000000000111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111100000000000011111111111111000000000000000000011111111111000000000000000000001111111", 
 "111111100000000000011111111111111000000000000000000011111111111000000000000000000001111111", 
 "111110000000000000000111111111100000000000000000000000111111100000000000000000000000111111", 
 "111100000001111000000111111111000000111111111111000000011111000000111111111111100000011111", 
 "111100000001111000000111111111000000111111111111100000011111000000111111111111100000011111", 
 "111100001111111000000111111111000000111000000011100000000111000000111000000001100000000111", 
 "111100001111111000000111111111000111110000000001111100000111000011111000000001111100000011", 
 "111100000011111000000111111111000111110000000001111100000111000011111000000001111100000011", 
 "111100000001111000000111111111000111110000001111111100000111000011111000000111111100000011", 
 "111110000001111000000111111111000111110000001111111100000111000011111000001111111100000011", 
 "111111100001111000000111111111000111110000001111111100000111000011111000000111111100000011", 
 "111111100001111000000111111111000111110000110001111100000111000011111000110001111100000011", 
 "111111100001111000000111111111000111110000110001111100000111000011111000110001111100000011", 
 "111111100001111000000111111111000111110000000001111100000111000011111000000001111100000011", 
 "111111100001111000000111111111000111111110000001111100000111000011111110000001111100000011", 
 "110000000001111000000000111111000111111110000001111100000111000011111110000001111100000011", 
 "110000000001111000000000111111000111110000000001111100000111000011111000000001111100000011", 
 "110000000001111000000000111111000111110000000001111100000111000011111000000001111100000011", 
 "110000111111111111110000001111000011110000000001111000000111000011111000000001111100000011", 
 "110001111111111111111000000111000000111111111111100000000111000000111111111111100000000011", 
 "110001111111111111111000000111000000111111111111100000000111000000111111111111100000000011", 
 "110000000000000000000000000111000000100000000000000000000111000000100000000000000000000011", 
 "110000000000000000000000000111110000000000000000000000000111111000000000000000000000000011", 
 "110000000000000000000000000111111000000000000000000000000111111000000000000000000000000011", 
 "111100000000000000000000000111111000000000000000000000000111111100000000000000000000000111", 
 "111100000000000000000000000111111110000000000000000000011111111111000000000000000000011111", 
 "111111111111111111111111111111111110000000000000000000011111111111000000000000000000011111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111", 
 "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111");

zero_big <=
("11111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111000011110000000000000000000000000000001111000011111111111111111111",
 "11111111111100000000000000000000000000000000000000000000000001111111111111111111",
 "11111111111000000000000000000000000000000000000000000000000001111111111111111111",
 "11111111111000000000000000000000000000000000000000000000000001111111111111111111",
 "11111111111000000000000000000000000000000000000000000000000001111111111111111111",
 "11111111111000000000000000000000000000000000000000000000000000111111111111111111",
 "11111101000000000000000000000000000000000000000000000000000000000111111111111111",
 "11111000000000000000000000000000000000000000000000000000000000000000111111111111",
 "11111000000000000000000000000000000000000000000000000000000000000000011111111111",
 "11111000000000000000111111111111111111111111111111111000000000000000011111111111",
 "11111000000000000001111111111111111111111111111111111000000000000000011111111111",
 "11111000000000000001111111111111111111111111111111111000000000000000011111111111",
 "11111000000000000001111111111111111111111111111111111000000000000000011111111111",
 "11111000000000000001111111111111111111111111111111111000000000000000001111111111",
 "11111000000000000011111111000000000000000000000111111100000000000000000000111111",
 "11111000000001111111111111000000000000000000000011111111111100000000000000011111",
 "11111000000001111111111111000000000000000000000011111111111100000000000000011111",
 "11111000000001111111111111000000000000000000000011111111111100000000000000011111",
 "11111000000001111111111111000000000000000000000011111111111100000000000000011111",
 "11111000000001111111111111000000000000000000000111111111111100000000000000011111",
 "11111000000001111111111111000000000000000000000111111111111100000000000000011111",
 "11111000000001111111111111000000000000000000001111111111111100000000000000011111",
 "11111000000001111111111111000000000000000111111111111111111100000000000000011111",
 "11111000000001111111111111000000000000001111111111111111111100000000000000011111",
 "11111000000001111111111111000000000000001111111111111111111100000000000000011111",
 "11111000000001111111111111000000000000001111111111111111111100000000000000011111",
 "11111000000001111111111111000000000000001111111111111111111100000000000000011111",
 "11111000000001111111111111000000000000000100011111111111111100000000000000011111",
 "11111000000001111111111111000000000111100000000111111111111110000000000000011111",
 "11111000000001111111111111000000001111100000000011111111111100000000000000011111",
 "11111000000001111111111111000000001111100000000011111111111100000000000000011111",
 "11111000000001111111111111000000001111100000000011111111111100000000000000011111",
 "11111000000001111111111111000000001111100000000011111111111100000000000000011111",
 "11111000000001111111111111000000001111100000000011111111111100000000000000011111",
 "11111000000001111111111111000000000111100000000011111111111100000000000000011111",
 "11111000000001111111111111100000000000000000000011111111111100000000000000011111",
 "11111000000001111111111111111111000000000000000011111111111100000000000000011111",
 "11111000000001111111111111111111000000000000000011111111111100000000000000011111",
 "11111000000001111111111111111111000000000000000011111111111100000000000000011111",
 "11111000000001111111111111111111000000000000000011111111111100000000000000011111",
 "11111000000001111111111111111110000000000000000011111111111100000000000000011111",
 "11111000000001111111111111000000000000000000000011111111111100000000000000011111",
 "11111000000001111111111111000000000000000000000011111111111100000000000000011111",
 "11111000000001111111111111000000000000000000000011111111111100000000000000011111",
 "11111000000001111111111111000000000000000000000011111111111100000000000000011111",
 "11111000000001111111111111000000000000000000000011111111111100000000000000011111",
 "11111000000001111111111111000000000000000000000011111111111100000000000000011111",
 "11111000000001111111111111000000000000000000000011111111111100000000000000011111",
 "11111000000000000011111111000000000000000000000111111110000000000000000000011111",
 "11111000000000000001111111111111111111111111111111111100000000000000000000011111",
 "11111000000000000001111111111111111111111111111111111000000000000000000000011111",
 "11111000000000000001111111111111111111111111111111111000000000000000000000011111",
 "11111000000000000001111111111111111111111111111111111000000000000000000000011111",
 "11111000000000000001111111111111111111111111111111111000000000000000000000011111",
 "11111000000000000000111111111111111111111111111111111000000000000000000000011111",
 "11111000000000000000111111111111111111111111111111110000000000000000000000011111",
 "11111100000000000000000000000000000000000000000000000000000000000000000000011111",
 "11111111111000000000000000000000000000000000000000000000000000000000000000011111",
 "11111111111000000000000000000000000000000000000000000000000000000000000000011111",
 "11111111111000000000000000000000000000000000000000000000000000000000000000011111",
 "11111111111100000000000000000000000000000000000000000000000000000000000000011111",
 "11111111111100000000000000000000000000000000000000000000000000000000000000011111",
 "11111111111100000000000000000000000000000000000000000000000000000000000000111111",
 "11111111111111111000000000000000000000000000000000000000000000000000001111111111",
 "11111111111111111100000000000000000000000000000000000000000000000000011111111111",
 "11111111111111111110000000000000000000000000000000000000000000000000011111111111",
 "11111111111111111100000000000000000000000000000000000000000000000000011111111111",
 "11111111111111111110000000000000000000000000000000000000000000000000011111111111",
 "11111111111111111110000000000000000000000000000000000000000000000000011111111111",
 "11111111111111111110000000000000000000000000000000000000000000000000111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111");



One_big <=
("11111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111000000000000000000000000000011111111111111111111111111111",
 "11111111111111111111100000000000000000000000000000001111111111111111111111111111",
 "11111111111111111111100000000000000000000000000000001111111111111111111111111111",
 "11111111111111111111100000000000000000000000000000001111111111111111111111111111",
 "11111111111111111111100000000000000000000000000000001111111111111111111111111111",
 "11111111111111111111100000000000000000000000000000001111111111111111111111111111",
 "11111111111111111111000000000000000000000000000000000111111111111111111111111111",
 "11111111111111100000000000000000000000000000000000000000001111111111111111111111",
 "11111111111111000000000000000000000000000000000000000000001111111111111111111111",
 "11111111111111000000000000000001111111111100000000000000001111111111111111111111",
 "11111111111111000000000000000011111111111110000000000000001111111111111111111111",
 "11111111111111000000000000000011111111111110000000000000001111111111111111111111",
 "11111111111111000000000000000011111111111110000000000000001111111111111111111111",
 "11111111111111000000000000000011111111111110000000000000001111111111111111111111",
 "11111111111111000000000000000011111111111110000000000000001111111111111111111111",
 "11111111111111000000000000001111111111111110000000000000001111111111111111111111",
 "11111111111111000000001111111111111111111110000000000000001111111111111111111111",
 "11111111111111000000001111111111111111111110000000000000001111111111111111111111",
 "11111111111111000000001111111111111111111110000000000000001111111111111111111111",
 "11111111111111000000001111111111111111111110000000000000001111111111111111111111",
 "11111111111111000000000111111111111111111110000000000000001111111111111111111111",
 "11111111111111000000000000000111111111111110000000000000001111111111111111111111",
 "11111111111111000000000000000011111111111110000000000000001111111111111111111111",
 "11111111111111000000000000000011111111111110000000000000001111111111111111111111",
 "11111111111111000000000000000011111111111110000000000000001111111111111111111111",
 "11111111111111000000000000000011111111111110000000000000001111111111111111111111",
 "11111111111111000000000000000011111111111110000000000000001111111111111111111111",
 "11111111111111000000000000000011111111111110000000000000001111111111111111111111",
 "11111111111111000000000000000011111111111110000000000000001111111111111111111111",
 "11111111111111100000000000000011111111111110000000000000001111111111111111111111",
 "11111111111111111111100000000011111111111110000000000000001111111111111111111111",
 "11111111111111111111100000000011111111111110000000000000001111111111111111111111",
 "11111111111111111111100000000011111111111110000000000000001111111111111111111111",
 "11111111111111111111100000000011111111111110000000000000001111111111111111111111",
 "11111111111111111111100000000011111111111110000000000000001111111111111111111111",
 "11111111111111111111100000000011111111111110000000000000001111111111111111111111",
 "11111111111111111111100000000011111111111110000000000000001111111111111111111111",
 "11111111111111111111100000000011111111111110000000000000001111111111111111111111",
 "11111111111111111111100000000011111111111110000000000000001111111111111111111111",
 "11111111111111111111100000000011111111111110000000000000001111111111111111111111",
 "11111111111111111111100000000011111111111110000000000000001111111111111111111111",
 "11111111111111111111100000000011111111111110000000000000001111111111111111111111",
 "11111111111111111111100000000011111111111110000000000000000111111111111111111111",
 "11111111000000000000000000000011111111111110000000000000000000000111111111111111",
 "11111110000000000000000000000011111111111110000000000000000000000011111111111111",
 "11111110000000000000000000000011111111111110000000000000000000000011111111111111",
 "11111110000000000000000000000011111111111110000000000000000000000011111111111111",
 "11111110000000000000000000000011111111111110000000000000000000000001111111111111",
 "11111110000000000000000000000011111111111110000000000000000000000011111111111111",
 "11111110000000000000000000000011111111111110000000000000000000000011111111111111",
 "11111110000000000000000000000011111111111110000000000000000000000001111111111111",
 "11111110000000000000000000000011111111111110000000000000000000000000001111111111",
 "11111110000000000111111111111111111111111111111111111111100000000000000001111111",
 "11111110000000001111111111111111111111111111111111111111110000000000000000111111",
 "11111110000000001111111111111111111111111111111111111111110000000000000000111111",
 "11111110000000001111111111111111111111111111111111111111100000000000000000111111",
 "11111110000000001111111111111111111111111111111111111111100000000000000000111111",
 "11111110000000001111111111111111111111111111111111111111100000000000000000111111",
 "11111110000000001111111111111111111111111111111111111111100000000000000000111111",
 "11111110000000000000000000000000000000000000000000000000000000000000000000111111",
 "11111110000000000000000000000000000000000000000000000000000000000000000000111111",
 "11111110000000000000000000000000000000000000000000000000000000000000000000111111",
 "11111110000000000000000000000000000000000000000000000000000000000000000000111111",
 "11111110000000000000000000000000000000000000000000000000000000000000000000111111",
 "11111110000000000000000000000000000000000000000000000000000000000000000000111111",
 "11111110000000000000000000000000000000000000000000000000000000000000000000111111",
 "11111110000000000000000000000000000000000000000000000000000000000000000000111111",
 "11111111000000000000000000000000000000000000000000000000000000000000000000111111",
 "11111111111110000000000000000000000000000000000000000000000000000000000000111111",
 "11111111111111000000000000000000000000000000000000000000000000000000000000111111",
 "11111111111111000000000000000000000000000000000000000000000000000000000000111111",
 "11111111111111000000000000000000000000000000000000000000000000000000000000111111",
 "11111111111111000000000000000000000000000000000000000000000000000000000000111111",
 "11111111111111000000000000000000000000000000000000000000000000000000000000111111",
 "11111111111111110000000000000000000000000000000000000000000000000000000011111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111",
 "11111111111111111111111111111111111111111111111111111111111111111111111111111111");

end Behavioral;                                                                                                                                                                                           
                                                                                                                                                                                                             
                                                                                                                                                                                                             